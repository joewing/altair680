

module basic_rom(addr_in, data_out);

   input wire [12:0] addr_in;
   output reg [7:0] data_out;

   always @(*) begin
      case (addr_in)
         0: data_out <= 8'h0d;
         1: data_out <= 8'h76;
         2: data_out <= 8'h00;
         3: data_out <= 8'hf3;
         4: data_out <= 8'h7e;
         5: data_out <= 8'h1a;
         6: data_out <= 8'h4f;
         7: data_out <= 8'h7e;
         8: data_out <= 8'h03;
         9: data_out <= 8'h4a;
         10: data_out <= 8'h00;
         11: data_out <= 8'h00;
         12: data_out <= 8'h48;
         13: data_out <= 8'h38;
         14: data_out <= 8'h00;
         15: data_out <= 8'h2c;
         16: data_out <= 8'h00;
         17: data_out <= 8'h00;
         18: data_out <= 8'h00;
         19: data_out <= 8'h00;
         20: data_out <= 8'h00;
         21: data_out <= 8'h00;
         22: data_out <= 8'h00;
         23: data_out <= 8'h00;
         24: data_out <= 8'h00;
         25: data_out <= 8'h00;
         26: data_out <= 8'h00;
         27: data_out <= 8'h00;
         28: data_out <= 8'h00;
         29: data_out <= 8'h00;
         30: data_out <= 8'h00;
         31: data_out <= 8'h00;
         32: data_out <= 8'h00;
         33: data_out <= 8'h00;
         34: data_out <= 8'h00;
         35: data_out <= 8'h00;
         36: data_out <= 8'h00;
         37: data_out <= 8'h00;
         38: data_out <= 8'h00;
         39: data_out <= 8'h00;
         40: data_out <= 8'h00;
         41: data_out <= 8'h00;
         42: data_out <= 8'h00;
         43: data_out <= 8'h00;
         44: data_out <= 8'h00;
         45: data_out <= 8'h00;
         46: data_out <= 8'h00;
         47: data_out <= 8'h00;
         48: data_out <= 8'h00;
         49: data_out <= 8'h00;
         50: data_out <= 8'h00;
         51: data_out <= 8'h00;
         52: data_out <= 8'h00;
         53: data_out <= 8'h00;
         54: data_out <= 8'h00;
         55: data_out <= 8'h00;
         56: data_out <= 8'h00;
         57: data_out <= 8'h00;
         58: data_out <= 8'h00;
         59: data_out <= 8'h00;
         60: data_out <= 8'h00;
         61: data_out <= 8'h00;
         62: data_out <= 8'h00;
         63: data_out <= 8'h00;
         64: data_out <= 8'h00;
         65: data_out <= 8'h00;
         66: data_out <= 8'h00;
         67: data_out <= 8'h00;
         68: data_out <= 8'h00;
         69: data_out <= 8'h00;
         70: data_out <= 8'h00;
         71: data_out <= 8'h00;
         72: data_out <= 8'h00;
         73: data_out <= 8'h00;
         74: data_out <= 8'h00;
         75: data_out <= 8'h00;
         76: data_out <= 8'h00;
         77: data_out <= 8'h00;
         78: data_out <= 8'h00;
         79: data_out <= 8'h00;
         80: data_out <= 8'h00;
         81: data_out <= 8'h00;
         82: data_out <= 8'h00;
         83: data_out <= 8'h00;
         84: data_out <= 8'h00;
         85: data_out <= 8'h00;
         86: data_out <= 8'h00;
         87: data_out <= 8'h00;
         88: data_out <= 8'h00;
         89: data_out <= 8'h00;
         90: data_out <= 8'h00;
         91: data_out <= 8'h00;
         92: data_out <= 8'h00;
         93: data_out <= 8'h00;
         94: data_out <= 8'h00;
         95: data_out <= 8'h00;
         96: data_out <= 8'h00;
         97: data_out <= 8'h00;
         98: data_out <= 8'h00;
         99: data_out <= 8'h00;
         100: data_out <= 8'h00;
         101: data_out <= 8'h00;
         102: data_out <= 8'h00;
         103: data_out <= 8'h00;
         104: data_out <= 8'h00;
         105: data_out <= 8'h00;
         106: data_out <= 8'h00;
         107: data_out <= 8'h00;
         108: data_out <= 8'h00;
         109: data_out <= 8'h00;
         110: data_out <= 8'h00;
         111: data_out <= 8'h00;
         112: data_out <= 8'h00;
         113: data_out <= 8'h00;
         114: data_out <= 8'h00;
         115: data_out <= 8'h00;
         116: data_out <= 8'h00;
         117: data_out <= 8'h00;
         118: data_out <= 8'h00;
         119: data_out <= 8'h00;
         120: data_out <= 8'h00;
         121: data_out <= 8'h00;
         122: data_out <= 8'h00;
         123: data_out <= 8'h00;
         124: data_out <= 8'h00;
         125: data_out <= 8'h00;
         126: data_out <= 8'h00;
         127: data_out <= 8'h00;
         128: data_out <= 8'h00;
         129: data_out <= 8'h00;
         130: data_out <= 8'h00;
         131: data_out <= 8'h00;
         132: data_out <= 8'h00;
         133: data_out <= 8'h00;
         134: data_out <= 8'h00;
         135: data_out <= 8'h00;
         136: data_out <= 8'h00;
         137: data_out <= 8'h00;
         138: data_out <= 8'h00;
         139: data_out <= 8'h00;
         140: data_out <= 8'h00;
         141: data_out <= 8'h00;
         142: data_out <= 8'h00;
         143: data_out <= 8'h00;
         144: data_out <= 8'h00;
         145: data_out <= 8'h00;
         146: data_out <= 8'h00;
         147: data_out <= 8'h00;
         148: data_out <= 8'h00;
         149: data_out <= 8'h00;
         150: data_out <= 8'h00;
         151: data_out <= 8'h00;
         152: data_out <= 8'h00;
         153: data_out <= 8'h00;
         154: data_out <= 8'h00;
         155: data_out <= 8'h00;
         156: data_out <= 8'h00;
         157: data_out <= 8'h00;
         158: data_out <= 8'h00;
         159: data_out <= 8'h00;
         160: data_out <= 8'h00;
         161: data_out <= 8'h00;
         162: data_out <= 8'h00;
         163: data_out <= 8'h00;
         164: data_out <= 8'h00;
         165: data_out <= 8'h00;
         166: data_out <= 8'h00;
         167: data_out <= 8'h00;
         168: data_out <= 8'h00;
         169: data_out <= 8'h00;
         170: data_out <= 8'h00;
         171: data_out <= 8'h00;
         172: data_out <= 8'h00;
         173: data_out <= 8'h00;
         174: data_out <= 8'h00;
         175: data_out <= 8'h00;
         176: data_out <= 8'h00;
         177: data_out <= 8'h00;
         178: data_out <= 8'h00;
         179: data_out <= 8'h00;
         180: data_out <= 8'h00;
         181: data_out <= 8'h00;
         182: data_out <= 8'h00;
         183: data_out <= 8'h00;
         184: data_out <= 8'h00;
         185: data_out <= 8'h00;
         186: data_out <= 8'h00;
         187: data_out <= 8'h00;
         188: data_out <= 8'h00;
         189: data_out <= 8'h00;
         190: data_out <= 8'h00;
         191: data_out <= 8'h7c;
         192: data_out <= 8'h00;
         193: data_out <= 8'hc9;
         194: data_out <= 8'h26;
         195: data_out <= 8'h03;
         196: data_out <= 8'h7c;
         197: data_out <= 8'h00;
         198: data_out <= 8'hc8;
         199: data_out <= 8'hb6;
         200: data_out <= 8'hea;
         201: data_out <= 8'h60;
         202: data_out <= 8'h81;
         203: data_out <= 8'h3a;
         204: data_out <= 8'h24;
         205: data_out <= 8'h08;
         206: data_out <= 8'h81;
         207: data_out <= 8'h20;
         208: data_out <= 8'h27;
         209: data_out <= 8'hed;
         210: data_out <= 8'h80;
         211: data_out <= 8'h30;
         212: data_out <= 8'h80;
         213: data_out <= 8'hd0;
         214: data_out <= 8'h39;
         215: data_out <= 8'hff;
         216: data_out <= 8'hea;
         217: data_out <= 8'h60;
         218: data_out <= 8'h7e;
         219: data_out <= 8'h03;
         220: data_out <= 8'hd5;
         221: data_out <= 8'h00;
         222: data_out <= 8'h00;
         223: data_out <= 8'h00;
         224: data_out <= 8'h00;
         225: data_out <= 8'h00;
         226: data_out <= 8'h00;
         227: data_out <= 8'h00;
         228: data_out <= 8'h00;
         229: data_out <= 8'h00;
         230: data_out <= 8'h00;
         231: data_out <= 8'h00;
         232: data_out <= 8'h00;
         233: data_out <= 8'h00;
         234: data_out <= 8'h00;
         235: data_out <= 8'h00;
         236: data_out <= 8'h00;
         237: data_out <= 8'h00;
         238: data_out <= 8'h00;
         239: data_out <= 8'h00;
         240: data_out <= 8'h00;
         241: data_out <= 8'h00;
         242: data_out <= 8'h00;
         243: data_out <= 8'h00;
         244: data_out <= 8'h00;
         245: data_out <= 8'h00;
         246: data_out <= 8'h00;
         247: data_out <= 8'h00;
         248: data_out <= 8'h00;
         249: data_out <= 8'h00;
         250: data_out <= 8'h00;
         251: data_out <= 8'h00;
         252: data_out <= 8'h00;
         253: data_out <= 8'h00;
         254: data_out <= 8'h00;
         255: data_out <= 8'h00;
         256: data_out <= 8'h00;
         257: data_out <= 8'h00;
         258: data_out <= 8'h00;
         259: data_out <= 8'h00;
         260: data_out <= 8'h00;
         261: data_out <= 8'h00;
         262: data_out <= 8'h00;
         263: data_out <= 8'h00;
         264: data_out <= 8'h00;
         265: data_out <= 8'h00;
         266: data_out <= 8'h00;
         267: data_out <= 8'h00;
         268: data_out <= 8'h00;
         269: data_out <= 8'h80;
         270: data_out <= 8'h4f;
         271: data_out <= 8'hc7;
         272: data_out <= 8'h52;
         273: data_out <= 8'h00;
         274: data_out <= 8'h7e;
         275: data_out <= 8'h1a;
         276: data_out <= 8'h4f;
         277: data_out <= 8'h0c;
         278: data_out <= 8'hf1;
         279: data_out <= 8'h0e;
         280: data_out <= 8'h60;
         281: data_out <= 8'h15;
         282: data_out <= 8'he6;
         283: data_out <= 8'h16;
         284: data_out <= 8'h5a;
         285: data_out <= 8'h16;
         286: data_out <= 8'h00;
         287: data_out <= 8'h0d;
         288: data_out <= 8'h71;
         289: data_out <= 8'h0e;
         290: data_out <= 8'h41;
         291: data_out <= 8'h0e;
         292: data_out <= 8'h6c;
         293: data_out <= 8'h18;
         294: data_out <= 8'h52;
         295: data_out <= 8'h19;
         296: data_out <= 8'h32;
         297: data_out <= 8'h14;
         298: data_out <= 8'h28;
         299: data_out <= 8'h18;
         300: data_out <= 8'hbe;
         301: data_out <= 8'h19;
         302: data_out <= 8'h68;
         303: data_out <= 8'h19;
         304: data_out <= 8'h6e;
         305: data_out <= 8'h19;
         306: data_out <= 8'hb4;
         307: data_out <= 8'h19;
         308: data_out <= 8'hf8;
         309: data_out <= 8'h11;
         310: data_out <= 8'hbc;
         311: data_out <= 8'h10;
         312: data_out <= 8'hd5;
         313: data_out <= 8'h0f;
         314: data_out <= 8'h1d;
         315: data_out <= 8'h11;
         316: data_out <= 8'h79;
         317: data_out <= 8'h10;
         318: data_out <= 8'hf5;
         319: data_out <= 8'h10;
         320: data_out <= 8'he1;
         321: data_out <= 8'h11;
         322: data_out <= 8'h00;
         323: data_out <= 8'h11;
         324: data_out <= 8'h1d;
         325: data_out <= 8'h11;
         326: data_out <= 8'h24;
         327: data_out <= 8'h79;
         328: data_out <= 8'h13;
         329: data_out <= 8'h1d;
         330: data_out <= 8'h79;
         331: data_out <= 8'h13;
         332: data_out <= 8'h12;
         333: data_out <= 8'h7b;
         334: data_out <= 8'h14;
         335: data_out <= 8'h60;
         336: data_out <= 8'h7b;
         337: data_out <= 8'h15;
         338: data_out <= 8'h14;
         339: data_out <= 8'h7f;
         340: data_out <= 8'h18;
         341: data_out <= 8'h5b;
         342: data_out <= 8'h50;
         343: data_out <= 8'h0b;
         344: data_out <= 8'ha4;
         345: data_out <= 8'h46;
         346: data_out <= 8'h0b;
         347: data_out <= 8'ha3;
         348: data_out <= 8'h45;
         349: data_out <= 8'h4e;
         350: data_out <= 8'hc4;
         351: data_out <= 8'h46;
         352: data_out <= 8'h4f;
         353: data_out <= 8'hd2;
         354: data_out <= 8'h4e;
         355: data_out <= 8'h45;
         356: data_out <= 8'h58;
         357: data_out <= 8'hd4;
         358: data_out <= 8'h44;
         359: data_out <= 8'h41;
         360: data_out <= 8'h54;
         361: data_out <= 8'hc1;
         362: data_out <= 8'h49;
         363: data_out <= 8'h4e;
         364: data_out <= 8'h50;
         365: data_out <= 8'h55;
         366: data_out <= 8'hd4;
         367: data_out <= 8'h44;
         368: data_out <= 8'h49;
         369: data_out <= 8'hcd;
         370: data_out <= 8'h52;
         371: data_out <= 8'h45;
         372: data_out <= 8'h41;
         373: data_out <= 8'hc4;
         374: data_out <= 8'h4c;
         375: data_out <= 8'h45;
         376: data_out <= 8'hd4;
         377: data_out <= 8'h47;
         378: data_out <= 8'h4f;
         379: data_out <= 8'h54;
         380: data_out <= 8'hcf;
         381: data_out <= 8'h52;
         382: data_out <= 8'h55;
         383: data_out <= 8'hce;
         384: data_out <= 8'h49;
         385: data_out <= 8'hc6;
         386: data_out <= 8'h52;
         387: data_out <= 8'h45;
         388: data_out <= 8'h53;
         389: data_out <= 8'h54;
         390: data_out <= 8'h4f;
         391: data_out <= 8'h52;
         392: data_out <= 8'hc5;
         393: data_out <= 8'h47;
         394: data_out <= 8'h4f;
         395: data_out <= 8'h53;
         396: data_out <= 8'h55;
         397: data_out <= 8'hc2;
         398: data_out <= 8'h52;
         399: data_out <= 8'h45;
         400: data_out <= 8'h54;
         401: data_out <= 8'h55;
         402: data_out <= 8'h52;
         403: data_out <= 8'hce;
         404: data_out <= 8'h52;
         405: data_out <= 8'h45;
         406: data_out <= 8'hcd;
         407: data_out <= 8'h53;
         408: data_out <= 8'h54;
         409: data_out <= 8'h4f;
         410: data_out <= 8'hd0;
         411: data_out <= 8'h4f;
         412: data_out <= 8'hce;
         413: data_out <= 8'h4e;
         414: data_out <= 8'h55;
         415: data_out <= 8'h4c;
         416: data_out <= 8'hcc;
         417: data_out <= 8'h57;
         418: data_out <= 8'h41;
         419: data_out <= 8'h49;
         420: data_out <= 8'hd4;
         421: data_out <= 8'h43;
         422: data_out <= 8'h4c;
         423: data_out <= 8'h4f;
         424: data_out <= 8'h41;
         425: data_out <= 8'hc4;
         426: data_out <= 8'h43;
         427: data_out <= 8'h53;
         428: data_out <= 8'h41;
         429: data_out <= 8'h56;
         430: data_out <= 8'hc5;
         431: data_out <= 8'h44;
         432: data_out <= 8'h45;
         433: data_out <= 8'hc6;
         434: data_out <= 8'h50;
         435: data_out <= 8'h4f;
         436: data_out <= 8'h4b;
         437: data_out <= 8'hc5;
         438: data_out <= 8'h50;
         439: data_out <= 8'h52;
         440: data_out <= 8'h49;
         441: data_out <= 8'h4e;
         442: data_out <= 8'hd4;
         443: data_out <= 8'h43;
         444: data_out <= 8'h4f;
         445: data_out <= 8'h4e;
         446: data_out <= 8'hd4;
         447: data_out <= 8'h4c;
         448: data_out <= 8'h49;
         449: data_out <= 8'h53;
         450: data_out <= 8'hd4;
         451: data_out <= 8'h43;
         452: data_out <= 8'h4c;
         453: data_out <= 8'h45;
         454: data_out <= 8'h41;
         455: data_out <= 8'hd2;
         456: data_out <= 8'h4e;
         457: data_out <= 8'h45;
         458: data_out <= 8'hd7;
         459: data_out <= 8'h54;
         460: data_out <= 8'h41;
         461: data_out <= 8'h42;
         462: data_out <= 8'ha8;
         463: data_out <= 8'h54;
         464: data_out <= 8'hcf;
         465: data_out <= 8'h46;
         466: data_out <= 8'hce;
         467: data_out <= 8'h53;
         468: data_out <= 8'h50;
         469: data_out <= 8'h43;
         470: data_out <= 8'ha8;
         471: data_out <= 8'h54;
         472: data_out <= 8'h48;
         473: data_out <= 8'h45;
         474: data_out <= 8'hce;
         475: data_out <= 8'h4e;
         476: data_out <= 8'h4f;
         477: data_out <= 8'hd4;
         478: data_out <= 8'h53;
         479: data_out <= 8'h54;
         480: data_out <= 8'h45;
         481: data_out <= 8'hd0;
         482: data_out <= 8'hab;
         483: data_out <= 8'had;
         484: data_out <= 8'haa;
         485: data_out <= 8'haf;
         486: data_out <= 8'hde;
         487: data_out <= 8'h41;
         488: data_out <= 8'h4e;
         489: data_out <= 8'hc4;
         490: data_out <= 8'h4f;
         491: data_out <= 8'hd2;
         492: data_out <= 8'hbe;
         493: data_out <= 8'hbd;
         494: data_out <= 8'hbc;
         495: data_out <= 8'h53;
         496: data_out <= 8'h47;
         497: data_out <= 8'hce;
         498: data_out <= 8'h49;
         499: data_out <= 8'h4e;
         500: data_out <= 8'hd4;
         501: data_out <= 8'h41;
         502: data_out <= 8'h42;
         503: data_out <= 8'hd3;
         504: data_out <= 8'h55;
         505: data_out <= 8'h53;
         506: data_out <= 8'hd2;
         507: data_out <= 8'h46;
         508: data_out <= 8'h52;
         509: data_out <= 8'hc5;
         510: data_out <= 8'h50;
         511: data_out <= 8'h4f;
         512: data_out <= 8'hd3;
         513: data_out <= 8'h53;
         514: data_out <= 8'h51;
         515: data_out <= 8'hd2;
         516: data_out <= 8'h52;
         517: data_out <= 8'h4e;
         518: data_out <= 8'hc4;
         519: data_out <= 8'h4c;
         520: data_out <= 8'h4f;
         521: data_out <= 8'hc7;
         522: data_out <= 8'h45;
         523: data_out <= 8'h58;
         524: data_out <= 8'hd0;
         525: data_out <= 8'h43;
         526: data_out <= 8'h4f;
         527: data_out <= 8'hd3;
         528: data_out <= 8'h53;
         529: data_out <= 8'h49;
         530: data_out <= 8'hce;
         531: data_out <= 8'h54;
         532: data_out <= 8'h41;
         533: data_out <= 8'hce;
         534: data_out <= 8'h41;
         535: data_out <= 8'h54;
         536: data_out <= 8'hce;
         537: data_out <= 8'h50;
         538: data_out <= 8'h45;
         539: data_out <= 8'h45;
         540: data_out <= 8'hcb;
         541: data_out <= 8'h4c;
         542: data_out <= 8'h45;
         543: data_out <= 8'hce;
         544: data_out <= 8'h53;
         545: data_out <= 8'h54;
         546: data_out <= 8'h52;
         547: data_out <= 8'ha4;
         548: data_out <= 8'h56;
         549: data_out <= 8'h41;
         550: data_out <= 8'hcc;
         551: data_out <= 8'h41;
         552: data_out <= 8'h53;
         553: data_out <= 8'hc3;
         554: data_out <= 8'h43;
         555: data_out <= 8'h48;
         556: data_out <= 8'h52;
         557: data_out <= 8'ha4;
         558: data_out <= 8'h4c;
         559: data_out <= 8'h45;
         560: data_out <= 8'h46;
         561: data_out <= 8'h54;
         562: data_out <= 8'ha4;
         563: data_out <= 8'h52;
         564: data_out <= 8'h49;
         565: data_out <= 8'h47;
         566: data_out <= 8'h48;
         567: data_out <= 8'h54;
         568: data_out <= 8'ha4;
         569: data_out <= 8'h4d;
         570: data_out <= 8'h49;
         571: data_out <= 8'h44;
         572: data_out <= 8'ha4;
         573: data_out <= 8'h00;
         574: data_out <= 8'h06;
         575: data_out <= 8'h3c;
         576: data_out <= 8'h05;
         577: data_out <= 8'h73;
         578: data_out <= 8'h09;
         579: data_out <= 8'hc1;
         580: data_out <= 8'h07;
         581: data_out <= 8'h14;
         582: data_out <= 8'h08;
         583: data_out <= 8'he8;
         584: data_out <= 8'h0c;
         585: data_out <= 8'h2e;
         586: data_out <= 8'h09;
         587: data_out <= 8'h0e;
         588: data_out <= 8'h07;
         589: data_out <= 8'h9f;
         590: data_out <= 8'h06;
         591: data_out <= 8'hd7;
         592: data_out <= 8'h06;
         593: data_out <= 8'hb1;
         594: data_out <= 8'h07;
         595: data_out <= 8'h35;
         596: data_out <= 8'h06;
         597: data_out <= 8'h20;
         598: data_out <= 8'h06;
         599: data_out <= 8'hbb;
         600: data_out <= 8'h06;
         601: data_out <= 8'hee;
         602: data_out <= 8'h07;
         603: data_out <= 8'h48;
         604: data_out <= 8'h06;
         605: data_out <= 8'h3b;
         606: data_out <= 8'h07;
         607: data_out <= 8'h55;
         608: data_out <= 8'h06;
         609: data_out <= 8'h72;
         610: data_out <= 8'h11;
         611: data_out <= 8'hca;
         612: data_out <= 8'h12;
         613: data_out <= 8'h06;
         614: data_out <= 8'h11;
         615: data_out <= 8'he3;
         616: data_out <= 8'h0e;
         617: data_out <= 8'h7b;
         618: data_out <= 8'h11;
         619: data_out <= 8'hc3;
         620: data_out <= 8'h08;
         621: data_out <= 8'h08;
         622: data_out <= 8'h06;
         623: data_out <= 8'h60;
         624: data_out <= 8'h05;
         625: data_out <= 8'h22;
         626: data_out <= 8'h06;
         627: data_out <= 8'h83;
         628: data_out <= 8'h04;
         629: data_out <= 8'hf0;
         630: data_out <= 8'h4e;
         631: data_out <= 8'hc6;
         632: data_out <= 8'h53;
         633: data_out <= 8'hce;
         634: data_out <= 8'h52;
         635: data_out <= 8'hc7;
         636: data_out <= 8'h4f;
         637: data_out <= 8'hc4;
         638: data_out <= 8'h46;
         639: data_out <= 8'hc3;
         640: data_out <= 8'h4f;
         641: data_out <= 8'hd6;
         642: data_out <= 8'h4f;
         643: data_out <= 8'hcd;
         644: data_out <= 8'h55;
         645: data_out <= 8'hd3;
         646: data_out <= 8'h42;
         647: data_out <= 8'hd3;
         648: data_out <= 8'h44;
         649: data_out <= 8'hc4;
         650: data_out <= 8'h2f;
         651: data_out <= 8'hb0;
         652: data_out <= 8'h49;
         653: data_out <= 8'hc4;
         654: data_out <= 8'h54;
         655: data_out <= 8'hcd;
         656: data_out <= 8'h4f;
         657: data_out <= 8'hd3;
         658: data_out <= 8'h4c;
         659: data_out <= 8'hd3;
         660: data_out <= 8'h53;
         661: data_out <= 8'hd4;
         662: data_out <= 8'h43;
         663: data_out <= 8'hce;
         664: data_out <= 8'h55;
         665: data_out <= 8'hc6;
         666: data_out <= 8'h20;
         667: data_out <= 8'h45;
         668: data_out <= 8'h52;
         669: data_out <= 8'h52;
         670: data_out <= 8'h4f;
         671: data_out <= 8'hd2;
         672: data_out <= 8'h00;
         673: data_out <= 8'h20;
         674: data_out <= 8'h49;
         675: data_out <= 8'h4e;
         676: data_out <= 8'ha0;
         677: data_out <= 8'h00;
         678: data_out <= 8'h0d;
         679: data_out <= 8'h0a;
         680: data_out <= 8'h4f;
         681: data_out <= 8'hcb;
         682: data_out <= 8'h0d;
         683: data_out <= 8'h0a;
         684: data_out <= 8'h00;
         685: data_out <= 8'h0d;
         686: data_out <= 8'h0a;
         687: data_out <= 8'h42;
         688: data_out <= 8'h52;
         689: data_out <= 8'h45;
         690: data_out <= 8'h41;
         691: data_out <= 8'hcb;
         692: data_out <= 8'h00;
         693: data_out <= 8'h30;
         694: data_out <= 8'h08;
         695: data_out <= 8'h08;
         696: data_out <= 8'h08;
         697: data_out <= 8'h08;
         698: data_out <= 8'hc6;
         699: data_out <= 8'h10;
         700: data_out <= 8'hdf;
         701: data_out <= 8'h71;
         702: data_out <= 8'ha6;
         703: data_out <= 8'h00;
         704: data_out <= 8'h80;
         705: data_out <= 8'h81;
         706: data_out <= 8'h26;
         707: data_out <= 8'h14;
         708: data_out <= 8'hee;
         709: data_out <= 8'h01;
         710: data_out <= 8'hdf;
         711: data_out <= 8'h73;
         712: data_out <= 8'hde;
         713: data_out <= 8'h9e;
         714: data_out <= 8'h27;
         715: data_out <= 8'h08;
         716: data_out <= 8'h9c;
         717: data_out <= 8'h73;
         718: data_out <= 8'h27;
         719: data_out <= 8'h08;
         720: data_out <= 8'h8d;
         721: data_out <= 8'h42;
         722: data_out <= 8'h20;
         723: data_out <= 8'he6;
         724: data_out <= 8'hde;
         725: data_out <= 8'h73;
         726: data_out <= 8'hdf;
         727: data_out <= 8'h9e;
         728: data_out <= 8'hde;
         729: data_out <= 8'h71;
         730: data_out <= 8'h4d;
         731: data_out <= 8'h39;
         732: data_out <= 8'h8d;
         733: data_out <= 8'h20;
         734: data_out <= 8'h07;
         735: data_out <= 8'h36;
         736: data_out <= 8'h9f;
         737: data_out <= 8'h78;
         738: data_out <= 8'h0f;
         739: data_out <= 8'h9e;
         740: data_out <= 8'ha3;
         741: data_out <= 8'hde;
         742: data_out <= 8'ha5;
         743: data_out <= 8'h08;
         744: data_out <= 8'h09;
         745: data_out <= 8'ha6;
         746: data_out <= 8'h00;
         747: data_out <= 8'h36;
         748: data_out <= 8'h9c;
         749: data_out <= 8'ha9;
         750: data_out <= 8'h26;
         751: data_out <= 8'hf8;
         752: data_out <= 8'h31;
         753: data_out <= 8'h9f;
         754: data_out <= 8'ha7;
         755: data_out <= 8'h9e;
         756: data_out <= 8'h78;
         757: data_out <= 8'h32;
         758: data_out <= 8'h06;
         759: data_out <= 8'h39;
         760: data_out <= 8'h4f;
         761: data_out <= 8'h58;
         762: data_out <= 8'hdb;
         763: data_out <= 8'h81;
         764: data_out <= 8'h99;
         765: data_out <= 8'h80;
         766: data_out <= 8'hcb;
         767: data_out <= 8'h26;
         768: data_out <= 8'h89;
         769: data_out <= 8'h00;
         770: data_out <= 8'h25;
         771: data_out <= 8'h1b;
         772: data_out <= 8'h9f;
         773: data_out <= 8'h78;
         774: data_out <= 8'h91;
         775: data_out <= 8'h78;
         776: data_out <= 8'h25;
         777: data_out <= 8'h06;
         778: data_out <= 8'h22;
         779: data_out <= 8'h13;
         780: data_out <= 8'hd1;
         781: data_out <= 8'h79;
         782: data_out <= 8'h22;
         783: data_out <= 8'h0f;
         784: data_out <= 8'h39;
         785: data_out <= 8'h4f;
         786: data_out <= 8'hdf;
         787: data_out <= 8'h71;
         788: data_out <= 8'hdb;
         789: data_out <= 8'h72;
         790: data_out <= 8'h99;
         791: data_out <= 8'h71;
         792: data_out <= 8'h97;
         793: data_out <= 8'h73;
         794: data_out <= 8'hd7;
         795: data_out <= 8'h74;
         796: data_out <= 8'hde;
         797: data_out <= 8'h73;
         798: data_out <= 8'h39;
         799: data_out <= 8'hc6;
         800: data_out <= 8'h0c;
         801: data_out <= 8'hbd;
         802: data_out <= 8'h05;
         803: data_out <= 8'h0e;
         804: data_out <= 8'h7f;
         805: data_out <= 8'h01;
         806: data_out <= 8'h11;
         807: data_out <= 8'hbd;
         808: data_out <= 8'h08;
         809: data_out <= 8'h42;
         810: data_out <= 8'hbd;
         811: data_out <= 8'h08;
         812: data_out <= 8'ha1;
         813: data_out <= 8'hce;
         814: data_out <= 8'h02;
         815: data_out <= 8'h76;
         816: data_out <= 8'h8d;
         817: data_out <= 8'hdf;
         818: data_out <= 8'ha6;
         819: data_out <= 8'h00;
         820: data_out <= 8'hbd;
         821: data_out <= 8'h08;
         822: data_out <= 8'ha3;
         823: data_out <= 8'ha6;
         824: data_out <= 8'h01;
         825: data_out <= 8'hbd;
         826: data_out <= 8'h08;
         827: data_out <= 8'ha3;
         828: data_out <= 8'hce;
         829: data_out <= 8'h02;
         830: data_out <= 8'h99;
         831: data_out <= 8'hbd;
         832: data_out <= 8'h08;
         833: data_out <= 8'h87;
         834: data_out <= 8'hde;
         835: data_out <= 8'h8a;
         836: data_out <= 8'h08;
         837: data_out <= 8'h27;
         838: data_out <= 8'h03;
         839: data_out <= 8'hbd;
         840: data_out <= 8'h17;
         841: data_out <= 8'h2d;
         842: data_out <= 8'h7f;
         843: data_out <= 8'h01;
         844: data_out <= 8'h11;
         845: data_out <= 8'hce;
         846: data_out <= 8'h02;
         847: data_out <= 8'ha5;
         848: data_out <= 8'hbd;
         849: data_out <= 8'h01;
         850: data_out <= 8'h12;
         851: data_out <= 8'h86;
         852: data_out <= 8'h2c;
         853: data_out <= 8'h97;
         854: data_out <= 8'h0f;
         855: data_out <= 8'hbd;
         856: data_out <= 8'h03;
         857: data_out <= 8'hfa;
         858: data_out <= 8'hdf;
         859: data_out <= 8'hc8;
         860: data_out <= 8'hbd;
         861: data_out <= 8'h00;
         862: data_out <= 8'hbf;
         863: data_out <= 8'h27;
         864: data_out <= 8'hf2;
         865: data_out <= 8'h25;
         866: data_out <= 8'h0b;
         867: data_out <= 8'hce;
         868: data_out <= 8'hff;
         869: data_out <= 8'hff;
         870: data_out <= 8'hdf;
         871: data_out <= 8'h8a;
         872: data_out <= 8'hbd;
         873: data_out <= 8'h04;
         874: data_out <= 8'h3c;
         875: data_out <= 8'h7e;
         876: data_out <= 8'h05;
         877: data_out <= 8'hfd;
         878: data_out <= 8'hbd;
         879: data_out <= 8'h07;
         880: data_out <= 8'h75;
         881: data_out <= 8'hde;
         882: data_out <= 8'h8e;
         883: data_out <= 8'hdf;
         884: data_out <= 8'h0e;
         885: data_out <= 8'hbd;
         886: data_out <= 8'h04;
         887: data_out <= 8'h3c;
         888: data_out <= 8'hd7;
         889: data_out <= 8'h5a;
         890: data_out <= 8'hbd;
         891: data_out <= 8'h04;
         892: data_out <= 8'hd2;
         893: data_out <= 8'h25;
         894: data_out <= 8'h22;
         895: data_out <= 8'hd6;
         896: data_out <= 8'haa;
         897: data_out <= 8'he0;
         898: data_out <= 8'h01;
         899: data_out <= 8'h86;
         900: data_out <= 8'hff;
         901: data_out <= 8'hdb;
         902: data_out <= 8'h7d;
         903: data_out <= 8'h99;
         904: data_out <= 8'h7c;
         905: data_out <= 8'h97;
         906: data_out <= 8'h7c;
         907: data_out <= 8'hd7;
         908: data_out <= 8'h7d;
         909: data_out <= 8'h07;
         910: data_out <= 8'h36;
         911: data_out <= 8'h9f;
         912: data_out <= 8'h78;
         913: data_out <= 8'h0f;
         914: data_out <= 8'hae;
         915: data_out <= 8'h00;
         916: data_out <= 8'h34;
         917: data_out <= 8'h32;
         918: data_out <= 8'ha7;
         919: data_out <= 8'h00;
         920: data_out <= 8'h08;
         921: data_out <= 8'h9c;
         922: data_out <= 8'h7c;
         923: data_out <= 8'h26;
         924: data_out <= 8'hf8;
         925: data_out <= 8'h9e;
         926: data_out <= 8'h78;
         927: data_out <= 8'h32;
         928: data_out <= 8'h06;
         929: data_out <= 8'h96;
         930: data_out <= 8'h10;
         931: data_out <= 8'h27;
         932: data_out <= 8'h2b;
         933: data_out <= 8'h96;
         934: data_out <= 8'h7c;
         935: data_out <= 8'hd6;
         936: data_out <= 8'h7d;
         937: data_out <= 8'h97;
         938: data_out <= 8'ha5;
         939: data_out <= 8'hd7;
         940: data_out <= 8'ha6;
         941: data_out <= 8'hdb;
         942: data_out <= 8'h5a;
         943: data_out <= 8'h89;
         944: data_out <= 8'h00;
         945: data_out <= 8'h97;
         946: data_out <= 8'ha3;
         947: data_out <= 8'hd7;
         948: data_out <= 8'ha4;
         949: data_out <= 8'hbd;
         950: data_out <= 8'h02;
         951: data_out <= 8'hdc;
         952: data_out <= 8'h07;
         953: data_out <= 8'h36;
         954: data_out <= 8'h9f;
         955: data_out <= 8'h78;
         956: data_out <= 8'h0f;
         957: data_out <= 8'h8e;
         958: data_out <= 8'h00;
         959: data_out <= 8'h0b;
         960: data_out <= 8'h32;
         961: data_out <= 8'ha7;
         962: data_out <= 8'h00;
         963: data_out <= 8'h08;
         964: data_out <= 8'h9c;
         965: data_out <= 8'ha7;
         966: data_out <= 8'h26;
         967: data_out <= 8'hf8;
         968: data_out <= 8'h9e;
         969: data_out <= 8'h78;
         970: data_out <= 8'h32;
         971: data_out <= 8'h07;
         972: data_out <= 8'hde;
         973: data_out <= 8'ha3;
         974: data_out <= 8'hdf;
         975: data_out <= 8'h7c;
         976: data_out <= 8'hbd;
         977: data_out <= 8'h04;
         978: data_out <= 8'hfc;
         979: data_out <= 8'hde;
         980: data_out <= 8'h7a;
         981: data_out <= 8'ha6;
         982: data_out <= 8'h00;
         983: data_out <= 8'haa;
         984: data_out <= 8'h01;
         985: data_out <= 8'h26;
         986: data_out <= 8'h03;
         987: data_out <= 8'h7e;
         988: data_out <= 8'h03;
         989: data_out <= 8'h53;
         990: data_out <= 8'hdf;
         991: data_out <= 8'hd8;
         992: data_out <= 8'h08;
         993: data_out <= 8'h08;
         994: data_out <= 8'h08;
         995: data_out <= 8'h08;
         996: data_out <= 8'h08;
         997: data_out <= 8'ha6;
         998: data_out <= 8'h00;
         999: data_out <= 8'h26;
         1000: data_out <= 8'hfb;
         1001: data_out <= 8'h08;
         1002: data_out <= 8'h7e;
         1003: data_out <= 8'h00;
         1004: data_out <= 8'hd7;
         1005: data_out <= 8'hbd;
         1006: data_out <= 8'h08;
         1007: data_out <= 8'ha3;
         1008: data_out <= 8'h09;
         1009: data_out <= 8'h5a;
         1010: data_out <= 8'h26;
         1011: data_out <= 8'h0b;
         1012: data_out <= 8'hbd;
         1013: data_out <= 8'h08;
         1014: data_out <= 8'ha3;
         1015: data_out <= 8'hbd;
         1016: data_out <= 8'h08;
         1017: data_out <= 8'h42;
         1018: data_out <= 8'hce;
         1019: data_out <= 8'h00;
         1020: data_out <= 8'h10;
         1021: data_out <= 8'hc6;
         1022: data_out <= 8'h01;
         1023: data_out <= 8'h8d;
         1024: data_out <= 8'h2b;
         1025: data_out <= 8'h81;
         1026: data_out <= 8'h07;
         1027: data_out <= 8'h27;
         1028: data_out <= 8'h14;
         1029: data_out <= 8'h81;
         1030: data_out <= 8'h0d;
         1031: data_out <= 8'h27;
         1032: data_out <= 8'h20;
         1033: data_out <= 8'h81;
         1034: data_out <= 8'h20;
         1035: data_out <= 8'h25;
         1036: data_out <= 8'hf2;
         1037: data_out <= 8'h81;
         1038: data_out <= 8'h7d;
         1039: data_out <= 8'h24;
         1040: data_out <= 8'hee;
         1041: data_out <= 8'h81;
         1042: data_out <= 8'h40;
         1043: data_out <= 8'h27;
         1044: data_out <= 8'hdf;
         1045: data_out <= 8'h81;
         1046: data_out <= 8'h5f;
         1047: data_out <= 8'h27;
         1048: data_out <= 8'hd4;
         1049: data_out <= 8'ha7;
         1050: data_out <= 8'h00;
         1051: data_out <= 8'hc1;
         1052: data_out <= 8'h48;
         1053: data_out <= 8'h24;
         1054: data_out <= 8'h03;
         1055: data_out <= 8'h08;
         1056: data_out <= 8'h5c;
         1057: data_out <= 8'h8c;
         1058: data_out <= 8'h86;
         1059: data_out <= 8'h07;
         1060: data_out <= 8'hbd;
         1061: data_out <= 8'h08;
         1062: data_out <= 8'ha3;
         1063: data_out <= 8'h20;
         1064: data_out <= 8'hd6;
         1065: data_out <= 8'h7e;
         1066: data_out <= 8'h08;
         1067: data_out <= 8'h3d;
         1068: data_out <= 8'h37;
         1069: data_out <= 8'hbd;
         1070: data_out <= 8'hff;
         1071: data_out <= 8'h00;
         1072: data_out <= 8'h17;
         1073: data_out <= 8'h33;
         1074: data_out <= 8'h84;
         1075: data_out <= 8'h7f;
         1076: data_out <= 8'h81;
         1077: data_out <= 8'h0f;
         1078: data_out <= 8'h26;
         1079: data_out <= 8'h03;
         1080: data_out <= 8'h73;
         1081: data_out <= 8'h01;
         1082: data_out <= 8'h11;
         1083: data_out <= 8'h39;
         1084: data_out <= 8'h7f;
         1085: data_out <= 8'h00;
         1086: data_out <= 8'h5d;
         1087: data_out <= 8'h7a;
         1088: data_out <= 8'h00;
         1089: data_out <= 8'hc9;
         1090: data_out <= 8'hce;
         1091: data_out <= 8'h00;
         1092: data_out <= 8'h0f;
         1093: data_out <= 8'hdf;
         1094: data_out <= 8'hbd;
         1095: data_out <= 8'h9f;
         1096: data_out <= 8'h78;
         1097: data_out <= 8'h07;
         1098: data_out <= 8'h97;
         1099: data_out <= 8'h5f;
         1100: data_out <= 8'h01;
         1101: data_out <= 8'h0f;
         1102: data_out <= 8'h9e;
         1103: data_out <= 8'hc8;
         1104: data_out <= 8'h33;
         1105: data_out <= 8'hc1;
         1106: data_out <= 8'h20;
         1107: data_out <= 8'h27;
         1108: data_out <= 8'h32;
         1109: data_out <= 8'hd7;
         1110: data_out <= 8'h59;
         1111: data_out <= 8'hc1;
         1112: data_out <= 8'h22;
         1113: data_out <= 8'h27;
         1114: data_out <= 8'h55;
         1115: data_out <= 8'h96;
         1116: data_out <= 8'h5d;
         1117: data_out <= 8'h26;
         1118: data_out <= 8'h28;
         1119: data_out <= 8'hc1;
         1120: data_out <= 8'h3f;
         1121: data_out <= 8'h26;
         1122: data_out <= 8'h04;
         1123: data_out <= 8'hc6;
         1124: data_out <= 8'h97;
         1125: data_out <= 8'h20;
         1126: data_out <= 8'h20;
         1127: data_out <= 8'hc1;
         1128: data_out <= 8'h30;
         1129: data_out <= 8'h25;
         1130: data_out <= 8'h04;
         1131: data_out <= 8'hc1;
         1132: data_out <= 8'h3c;
         1133: data_out <= 8'h25;
         1134: data_out <= 8'h18;
         1135: data_out <= 8'hce;
         1136: data_out <= 8'h01;
         1137: data_out <= 8'h5b;
         1138: data_out <= 8'h9e;
         1139: data_out <= 8'hc8;
         1140: data_out <= 8'h5f;
         1141: data_out <= 8'h08;
         1142: data_out <= 8'h32;
         1143: data_out <= 8'h81;
         1144: data_out <= 8'h20;
         1145: data_out <= 8'h27;
         1146: data_out <= 8'hfb;
         1147: data_out <= 8'ha0;
         1148: data_out <= 8'h00;
         1149: data_out <= 8'h27;
         1150: data_out <= 8'hf6;
         1151: data_out <= 8'h81;
         1152: data_out <= 8'h80;
         1153: data_out <= 8'h26;
         1154: data_out <= 8'h32;
         1155: data_out <= 8'hca;
         1156: data_out <= 8'h80;
         1157: data_out <= 8'hde;
         1158: data_out <= 8'hbd;
         1159: data_out <= 8'h9f;
         1160: data_out <= 8'hc8;
         1161: data_out <= 8'h9e;
         1162: data_out <= 8'h78;
         1163: data_out <= 8'h96;
         1164: data_out <= 8'h5f;
         1165: data_out <= 8'h06;
         1166: data_out <= 8'h08;
         1167: data_out <= 8'hdf;
         1168: data_out <= 8'hbd;
         1169: data_out <= 8'he7;
         1170: data_out <= 8'h00;
         1171: data_out <= 8'h27;
         1172: data_out <= 8'h2f;
         1173: data_out <= 8'hc0;
         1174: data_out <= 8'h3a;
         1175: data_out <= 8'h27;
         1176: data_out <= 8'h04;
         1177: data_out <= 8'hc1;
         1178: data_out <= 8'h49;
         1179: data_out <= 8'h26;
         1180: data_out <= 8'h02;
         1181: data_out <= 8'hd7;
         1182: data_out <= 8'h5d;
         1183: data_out <= 8'hc0;
         1184: data_out <= 8'h54;
         1185: data_out <= 8'h26;
         1186: data_out <= 8'ha9;
         1187: data_out <= 8'hd7;
         1188: data_out <= 8'h59;
         1189: data_out <= 8'h0f;
         1190: data_out <= 8'h9e;
         1191: data_out <= 8'hc8;
         1192: data_out <= 8'h33;
         1193: data_out <= 8'h5d;
         1194: data_out <= 8'h27;
         1195: data_out <= 8'hdb;
         1196: data_out <= 8'hd1;
         1197: data_out <= 8'h59;
         1198: data_out <= 8'h27;
         1199: data_out <= 8'hd7;
         1200: data_out <= 8'h08;
         1201: data_out <= 8'he7;
         1202: data_out <= 8'h00;
         1203: data_out <= 8'h20;
         1204: data_out <= 8'hf3;
         1205: data_out <= 8'h9e;
         1206: data_out <= 8'hc8;
         1207: data_out <= 8'h5c;
         1208: data_out <= 8'ha6;
         1209: data_out <= 8'h00;
         1210: data_out <= 8'h08;
         1211: data_out <= 8'h2a;
         1212: data_out <= 8'hfb;
         1213: data_out <= 8'ha6;
         1214: data_out <= 8'h00;
         1215: data_out <= 8'h26;
         1216: data_out <= 8'hb5;
         1217: data_out <= 8'h33;
         1218: data_out <= 8'h20;
         1219: data_out <= 8'hc1;
         1220: data_out <= 8'he7;
         1221: data_out <= 8'h01;
         1222: data_out <= 8'he7;
         1223: data_out <= 8'h02;
         1224: data_out <= 8'hd6;
         1225: data_out <= 8'hbe;
         1226: data_out <= 8'hc0;
         1227: data_out <= 8'h0b;
         1228: data_out <= 8'hce;
         1229: data_out <= 8'h00;
         1230: data_out <= 8'h0f;
         1231: data_out <= 8'hdf;
         1232: data_out <= 8'hc8;
         1233: data_out <= 8'h39;
         1234: data_out <= 8'h96;
         1235: data_out <= 8'h8e;
         1236: data_out <= 8'hde;
         1237: data_out <= 8'h7a;
         1238: data_out <= 8'he6;
         1239: data_out <= 8'h00;
         1240: data_out <= 8'hea;
         1241: data_out <= 8'h01;
         1242: data_out <= 8'h27;
         1243: data_out <= 8'h10;
         1244: data_out <= 8'ha1;
         1245: data_out <= 8'h02;
         1246: data_out <= 8'h22;
         1247: data_out <= 8'h08;
         1248: data_out <= 8'h25;
         1249: data_out <= 8'h0b;
         1250: data_out <= 8'hd6;
         1251: data_out <= 8'h8f;
         1252: data_out <= 8'he1;
         1253: data_out <= 8'h03;
         1254: data_out <= 8'h23;
         1255: data_out <= 8'h05;
         1256: data_out <= 8'hee;
         1257: data_out <= 8'h00;
         1258: data_out <= 8'h20;
         1259: data_out <= 8'hea;
         1260: data_out <= 8'h0d;
         1261: data_out <= 8'hdf;
         1262: data_out <= 8'ha9;
         1263: data_out <= 8'h39;
         1264: data_out <= 8'h26;
         1265: data_out <= 8'hfb;
         1266: data_out <= 8'hde;
         1267: data_out <= 8'h7a;
         1268: data_out <= 8'h6f;
         1269: data_out <= 8'h00;
         1270: data_out <= 8'h08;
         1271: data_out <= 8'h6f;
         1272: data_out <= 8'h00;
         1273: data_out <= 8'h08;
         1274: data_out <= 8'hdf;
         1275: data_out <= 8'h7c;
         1276: data_out <= 8'hde;
         1277: data_out <= 8'h7a;
         1278: data_out <= 8'h09;
         1279: data_out <= 8'hdf;
         1280: data_out <= 8'hc8;
         1281: data_out <= 8'hde;
         1282: data_out <= 8'h88;
         1283: data_out <= 8'hdf;
         1284: data_out <= 8'h84;
         1285: data_out <= 8'hbd;
         1286: data_out <= 8'h06;
         1287: data_out <= 8'h20;
         1288: data_out <= 8'hde;
         1289: data_out <= 8'h7c;
         1290: data_out <= 8'hdf;
         1291: data_out <= 8'h7e;
         1292: data_out <= 8'hdf;
         1293: data_out <= 8'h80;
         1294: data_out <= 8'hce;
         1295: data_out <= 8'h00;
         1296: data_out <= 8'h65;
         1297: data_out <= 8'hdf;
         1298: data_out <= 8'h61;
         1299: data_out <= 8'h30;
         1300: data_out <= 8'hee;
         1301: data_out <= 8'h00;
         1302: data_out <= 8'h9e;
         1303: data_out <= 8'h82;
         1304: data_out <= 8'h4f;
         1305: data_out <= 8'h36;
         1306: data_out <= 8'h97;
         1307: data_out <= 8'h90;
         1308: data_out <= 8'h97;
         1309: data_out <= 8'h91;
         1310: data_out <= 8'h97;
         1311: data_out <= 8'h5e;
         1312: data_out <= 8'h6e;
         1313: data_out <= 8'h00;
         1314: data_out <= 8'h22;
         1315: data_out <= 8'had;
         1316: data_out <= 8'hbd;
         1317: data_out <= 8'h07;
         1318: data_out <= 8'h75;
         1319: data_out <= 8'h26;
         1320: data_out <= 8'ha8;
         1321: data_out <= 8'h32;
         1322: data_out <= 8'h32;
         1323: data_out <= 8'h8d;
         1324: data_out <= 8'ha5;
         1325: data_out <= 8'ha6;
         1326: data_out <= 8'h00;
         1327: data_out <= 8'haa;
         1328: data_out <= 8'h01;
         1329: data_out <= 8'h26;
         1330: data_out <= 8'h03;
         1331: data_out <= 8'h7e;
         1332: data_out <= 8'h03;
         1333: data_out <= 8'h4a;
         1334: data_out <= 8'hbd;
         1335: data_out <= 8'h06;
         1336: data_out <= 8'h26;
         1337: data_out <= 8'hbd;
         1338: data_out <= 8'h08;
         1339: data_out <= 8'h42;
         1340: data_out <= 8'ha6;
         1341: data_out <= 8'h02;
         1342: data_out <= 8'he6;
         1343: data_out <= 8'h03;
         1344: data_out <= 8'h08;
         1345: data_out <= 8'h08;
         1346: data_out <= 8'h08;
         1347: data_out <= 8'h08;
         1348: data_out <= 8'hdf;
         1349: data_out <= 8'h71;
         1350: data_out <= 8'hbd;
         1351: data_out <= 8'h17;
         1352: data_out <= 8'h36;
         1353: data_out <= 8'h86;
         1354: data_out <= 8'h20;
         1355: data_out <= 8'hde;
         1356: data_out <= 8'h71;
         1357: data_out <= 8'hbd;
         1358: data_out <= 8'h08;
         1359: data_out <= 8'ha3;
         1360: data_out <= 8'ha6;
         1361: data_out <= 8'h00;
         1362: data_out <= 8'h08;
         1363: data_out <= 8'h4d;
         1364: data_out <= 8'h27;
         1365: data_out <= 8'hd7;
         1366: data_out <= 8'h2a;
         1367: data_out <= 8'hf5;
         1368: data_out <= 8'h80;
         1369: data_out <= 8'h7f;
         1370: data_out <= 8'hdf;
         1371: data_out <= 8'h71;
         1372: data_out <= 8'hce;
         1373: data_out <= 8'h01;
         1374: data_out <= 8'h5c;
         1375: data_out <= 8'h4a;
         1376: data_out <= 8'h27;
         1377: data_out <= 8'h07;
         1378: data_out <= 8'he6;
         1379: data_out <= 8'h00;
         1380: data_out <= 8'h08;
         1381: data_out <= 8'h2a;
         1382: data_out <= 8'hfb;
         1383: data_out <= 8'h20;
         1384: data_out <= 8'hf6;
         1385: data_out <= 8'ha6;
         1386: data_out <= 8'h00;
         1387: data_out <= 8'h2b;
         1388: data_out <= 8'hde;
         1389: data_out <= 8'h08;
         1390: data_out <= 8'hbd;
         1391: data_out <= 8'h08;
         1392: data_out <= 8'ha3;
         1393: data_out <= 8'h20;
         1394: data_out <= 8'hf6;
         1395: data_out <= 8'h86;
         1396: data_out <= 8'h80;
         1397: data_out <= 8'h97;
         1398: data_out <= 8'h5e;
         1399: data_out <= 8'hbd;
         1400: data_out <= 8'h07;
         1401: data_out <= 8'h9f;
         1402: data_out <= 8'hbd;
         1403: data_out <= 8'h02;
         1404: data_out <= 8'hb5;
         1405: data_out <= 8'h31;
         1406: data_out <= 8'h31;
         1407: data_out <= 8'h26;
         1408: data_out <= 8'h04;
         1409: data_out <= 8'hbd;
         1410: data_out <= 8'h03;
         1411: data_out <= 8'h14;
         1412: data_out <= 8'h35;
         1413: data_out <= 8'hc6;
         1414: data_out <= 8'h08;
         1415: data_out <= 8'hbd;
         1416: data_out <= 8'h02;
         1417: data_out <= 8'hf8;
         1418: data_out <= 8'hbd;
         1419: data_out <= 8'h07;
         1420: data_out <= 8'h19;
         1421: data_out <= 8'hdf;
         1422: data_out <= 8'h71;
         1423: data_out <= 8'hd6;
         1424: data_out <= 8'h72;
         1425: data_out <= 8'h37;
         1426: data_out <= 8'hd6;
         1427: data_out <= 8'h71;
         1428: data_out <= 8'h37;
         1429: data_out <= 8'hd6;
         1430: data_out <= 8'h8b;
         1431: data_out <= 8'h37;
         1432: data_out <= 8'hd6;
         1433: data_out <= 8'h8a;
         1434: data_out <= 8'h37;
         1435: data_out <= 8'hc6;
         1436: data_out <= 8'h9d;
         1437: data_out <= 8'hbd;
         1438: data_out <= 8'h0b;
         1439: data_out <= 8'h4d;
         1440: data_out <= 8'hbd;
         1441: data_out <= 8'h0a;
         1442: data_out <= 8'h1b;
         1443: data_out <= 8'hbd;
         1444: data_out <= 8'h0a;
         1445: data_out <= 8'h19;
         1446: data_out <= 8'hd6;
         1447: data_out <= 8'hb3;
         1448: data_out <= 8'hca;
         1449: data_out <= 8'h7f;
         1450: data_out <= 8'hd4;
         1451: data_out <= 8'hb0;
         1452: data_out <= 8'hd7;
         1453: data_out <= 8'hb0;
         1454: data_out <= 8'hce;
         1455: data_out <= 8'h05;
         1456: data_out <= 8'hb4;
         1457: data_out <= 8'h7e;
         1458: data_out <= 8'h0a;
         1459: data_out <= 8'hb9;
         1460: data_out <= 8'hce;
         1461: data_out <= 8'h14;
         1462: data_out <= 8'h07;
         1463: data_out <= 8'hbd;
         1464: data_out <= 8'h15;
         1465: data_out <= 8'h8e;
         1466: data_out <= 8'hbd;
         1467: data_out <= 8'h00;
         1468: data_out <= 8'hc7;
         1469: data_out <= 8'h81;
         1470: data_out <= 8'ha2;
         1471: data_out <= 8'h26;
         1472: data_out <= 8'h06;
         1473: data_out <= 8'hbd;
         1474: data_out <= 8'h00;
         1475: data_out <= 8'hbf;
         1476: data_out <= 8'hbd;
         1477: data_out <= 8'h0a;
         1478: data_out <= 8'h19;
         1479: data_out <= 8'hbd;
         1480: data_out <= 8'h15;
         1481: data_out <= 8'hd9;
         1482: data_out <= 8'hbd;
         1483: data_out <= 8'h0a;
         1484: data_out <= 8'hb3;
         1485: data_out <= 8'hd6;
         1486: data_out <= 8'h9f;
         1487: data_out <= 8'h37;
         1488: data_out <= 8'hd6;
         1489: data_out <= 8'h9e;
         1490: data_out <= 8'h37;
         1491: data_out <= 8'h86;
         1492: data_out <= 8'h81;
         1493: data_out <= 8'h36;
         1494: data_out <= 8'h8d;
         1495: data_out <= 8'h4e;
         1496: data_out <= 8'hde;
         1497: data_out <= 8'hc8;
         1498: data_out <= 8'hdf;
         1499: data_out <= 8'h92;
         1500: data_out <= 8'ha6;
         1501: data_out <= 8'h00;
         1502: data_out <= 8'h27;
         1503: data_out <= 8'h07;
         1504: data_out <= 8'h81;
         1505: data_out <= 8'h3a;
         1506: data_out <= 8'h27;
         1507: data_out <= 8'h19;
         1508: data_out <= 8'h7e;
         1509: data_out <= 8'h0b;
         1510: data_out <= 8'h57;
         1511: data_out <= 8'h08;
         1512: data_out <= 8'ha6;
         1513: data_out <= 8'h00;
         1514: data_out <= 8'h08;
         1515: data_out <= 8'haa;
         1516: data_out <= 8'h00;
         1517: data_out <= 8'h0c;
         1518: data_out <= 8'h07;
         1519: data_out <= 8'h27;
         1520: data_out <= 8'h54;
         1521: data_out <= 8'h08;
         1522: data_out <= 8'ha6;
         1523: data_out <= 8'h00;
         1524: data_out <= 8'h97;
         1525: data_out <= 8'h8a;
         1526: data_out <= 8'h08;
         1527: data_out <= 8'ha6;
         1528: data_out <= 8'h00;
         1529: data_out <= 8'h97;
         1530: data_out <= 8'h8b;
         1531: data_out <= 8'hdf;
         1532: data_out <= 8'hc8;
         1533: data_out <= 8'hbd;
         1534: data_out <= 8'h00;
         1535: data_out <= 8'hbf;
         1536: data_out <= 8'h8d;
         1537: data_out <= 8'h02;
         1538: data_out <= 8'h20;
         1539: data_out <= 8'hd2;
         1540: data_out <= 8'h27;
         1541: data_out <= 8'h6b;
         1542: data_out <= 8'h80;
         1543: data_out <= 8'h80;
         1544: data_out <= 8'h24;
         1545: data_out <= 8'h03;
         1546: data_out <= 8'h7e;
         1547: data_out <= 8'h07;
         1548: data_out <= 8'h9f;
         1549: data_out <= 8'h81;
         1550: data_out <= 8'h1c;
         1551: data_out <= 8'h24;
         1552: data_out <= 8'hd3;
         1553: data_out <= 8'h48;
         1554: data_out <= 8'h16;
         1555: data_out <= 8'hce;
         1556: data_out <= 8'h02;
         1557: data_out <= 8'h3e;
         1558: data_out <= 8'hbd;
         1559: data_out <= 8'h03;
         1560: data_out <= 8'h11;
         1561: data_out <= 8'hee;
         1562: data_out <= 8'h00;
         1563: data_out <= 8'hbd;
         1564: data_out <= 8'h00;
         1565: data_out <= 8'hbf;
         1566: data_out <= 8'h6e;
         1567: data_out <= 8'h00;
         1568: data_out <= 8'hde;
         1569: data_out <= 8'h7a;
         1570: data_out <= 8'h09;
         1571: data_out <= 8'hdf;
         1572: data_out <= 8'h96;
         1573: data_out <= 8'h39;
         1574: data_out <= 8'hbd;
         1575: data_out <= 8'hff;
         1576: data_out <= 8'h24;
         1577: data_out <= 8'h24;
         1578: data_out <= 8'hfa;
         1579: data_out <= 8'hbd;
         1580: data_out <= 8'h04;
         1581: data_out <= 8'h2c;
         1582: data_out <= 8'h36;
         1583: data_out <= 8'hb6;
         1584: data_out <= 8'hf0;
         1585: data_out <= 8'h02;
         1586: data_out <= 8'h84;
         1587: data_out <= 8'h02;
         1588: data_out <= 8'h32;
         1589: data_out <= 8'h27;
         1590: data_out <= 8'h02;
         1591: data_out <= 8'h86;
         1592: data_out <= 8'h03;
         1593: data_out <= 8'h81;
         1594: data_out <= 8'h03;
         1595: data_out <= 8'h0d;
         1596: data_out <= 8'h26;
         1597: data_out <= 8'h33;
         1598: data_out <= 8'h07;
         1599: data_out <= 8'hde;
         1600: data_out <= 8'hc8;
         1601: data_out <= 8'hdf;
         1602: data_out <= 8'h92;
         1603: data_out <= 8'h31;
         1604: data_out <= 8'h31;
         1605: data_out <= 8'hde;
         1606: data_out <= 8'h8a;
         1607: data_out <= 8'h08;
         1608: data_out <= 8'h27;
         1609: data_out <= 8'h07;
         1610: data_out <= 8'h09;
         1611: data_out <= 8'hdf;
         1612: data_out <= 8'h8c;
         1613: data_out <= 8'hde;
         1614: data_out <= 8'h92;
         1615: data_out <= 8'hdf;
         1616: data_out <= 8'h90;
         1617: data_out <= 8'h7f;
         1618: data_out <= 8'h01;
         1619: data_out <= 8'h11;
         1620: data_out <= 8'hce;
         1621: data_out <= 8'h02;
         1622: data_out <= 8'hac;
         1623: data_out <= 8'h06;
         1624: data_out <= 8'h24;
         1625: data_out <= 8'h03;
         1626: data_out <= 8'h7e;
         1627: data_out <= 8'h03;
         1628: data_out <= 8'h3f;
         1629: data_out <= 8'h7e;
         1630: data_out <= 8'h03;
         1631: data_out <= 8'h4a;
         1632: data_out <= 8'h26;
         1633: data_out <= 8'h0f;
         1634: data_out <= 8'hc6;
         1635: data_out <= 8'h20;
         1636: data_out <= 8'hde;
         1637: data_out <= 8'h90;
         1638: data_out <= 8'h26;
         1639: data_out <= 8'h03;
         1640: data_out <= 8'h7e;
         1641: data_out <= 8'h03;
         1642: data_out <= 8'h21;
         1643: data_out <= 8'hdf;
         1644: data_out <= 8'hc8;
         1645: data_out <= 8'hde;
         1646: data_out <= 8'h8c;
         1647: data_out <= 8'hdf;
         1648: data_out <= 8'h8a;
         1649: data_out <= 8'h39;
         1650: data_out <= 8'hbd;
         1651: data_out <= 8'h11;
         1652: data_out <= 8'h6a;
         1653: data_out <= 8'h26;
         1654: data_out <= 8'hfa;
         1655: data_out <= 8'h5c;
         1656: data_out <= 8'hd1;
         1657: data_out <= 8'h0c;
         1658: data_out <= 8'h24;
         1659: data_out <= 8'h04;
         1660: data_out <= 8'h5a;
         1661: data_out <= 8'hd7;
         1662: data_out <= 8'h0a;
         1663: data_out <= 8'h39;
         1664: data_out <= 8'h7e;
         1665: data_out <= 8'h0d;
         1666: data_out <= 8'h71;
         1667: data_out <= 8'h27;
         1668: data_out <= 8'h29;
         1669: data_out <= 8'hbd;
         1670: data_out <= 8'h0c;
         1671: data_out <= 8'he7;
         1672: data_out <= 8'hbd;
         1673: data_out <= 8'h00;
         1674: data_out <= 8'hc7;
         1675: data_out <= 8'h26;
         1676: data_out <= 8'he4;
         1677: data_out <= 8'h96;
         1678: data_out <= 8'h88;
         1679: data_out <= 8'hd6;
         1680: data_out <= 8'h89;
         1681: data_out <= 8'hd0;
         1682: data_out <= 8'hb2;
         1683: data_out <= 8'h92;
         1684: data_out <= 8'hb1;
         1685: data_out <= 8'h25;
         1686: data_out <= 8'h14;
         1687: data_out <= 8'hde;
         1688: data_out <= 8'h82;
         1689: data_out <= 8'h97;
         1690: data_out <= 8'h82;
         1691: data_out <= 8'hd7;
         1692: data_out <= 8'h83;
         1693: data_out <= 8'hc0;
         1694: data_out <= 8'h28;
         1695: data_out <= 8'h82;
         1696: data_out <= 8'h00;
         1697: data_out <= 8'h25;
         1698: data_out <= 8'h06;
         1699: data_out <= 8'hd0;
         1700: data_out <= 8'h7d;
         1701: data_out <= 8'h92;
         1702: data_out <= 8'h7c;
         1703: data_out <= 8'h24;
         1704: data_out <= 8'h05;
         1705: data_out <= 8'hdf;
         1706: data_out <= 8'h82;
         1707: data_out <= 8'h7e;
         1708: data_out <= 8'h03;
         1709: data_out <= 8'h1f;
         1710: data_out <= 8'h7e;
         1711: data_out <= 8'h05;
         1712: data_out <= 8'h01;
         1713: data_out <= 8'h26;
         1714: data_out <= 8'h03;
         1715: data_out <= 8'h7e;
         1716: data_out <= 8'h04;
         1717: data_out <= 8'hfc;
         1718: data_out <= 8'hbd;
         1719: data_out <= 8'h05;
         1720: data_out <= 8'h01;
         1721: data_out <= 8'h20;
         1722: data_out <= 8'h14;
         1723: data_out <= 8'hc6;
         1724: data_out <= 8'h03;
         1725: data_out <= 8'hbd;
         1726: data_out <= 8'h02;
         1727: data_out <= 8'hf8;
         1728: data_out <= 8'hd6;
         1729: data_out <= 8'hc9;
         1730: data_out <= 8'h37;
         1731: data_out <= 8'hd6;
         1732: data_out <= 8'hc8;
         1733: data_out <= 8'h37;
         1734: data_out <= 8'hd6;
         1735: data_out <= 8'h8b;
         1736: data_out <= 8'h37;
         1737: data_out <= 8'hd6;
         1738: data_out <= 8'h8a;
         1739: data_out <= 8'h37;
         1740: data_out <= 8'h86;
         1741: data_out <= 8'h8c;
         1742: data_out <= 8'h36;
         1743: data_out <= 8'hbd;
         1744: data_out <= 8'h00;
         1745: data_out <= 8'hc7;
         1746: data_out <= 8'h8d;
         1747: data_out <= 8'h03;
         1748: data_out <= 8'h7e;
         1749: data_out <= 8'h05;
         1750: data_out <= 8'hd6;
         1751: data_out <= 8'hbd;
         1752: data_out <= 8'h07;
         1753: data_out <= 8'h75;
         1754: data_out <= 8'h8d;
         1755: data_out <= 8'h40;
         1756: data_out <= 8'h08;
         1757: data_out <= 8'h96;
         1758: data_out <= 8'h8e;
         1759: data_out <= 8'h91;
         1760: data_out <= 8'h8a;
         1761: data_out <= 8'h22;
         1762: data_out <= 8'h02;
         1763: data_out <= 8'hde;
         1764: data_out <= 8'h7a;
         1765: data_out <= 8'hbd;
         1766: data_out <= 8'h04;
         1767: data_out <= 8'hd6;
         1768: data_out <= 8'h25;
         1769: data_out <= 8'h15;
         1770: data_out <= 8'h09;
         1771: data_out <= 8'hdf;
         1772: data_out <= 8'hc8;
         1773: data_out <= 8'h39;
         1774: data_out <= 8'h26;
         1775: data_out <= 8'hfd;
         1776: data_out <= 8'h86;
         1777: data_out <= 8'hff;
         1778: data_out <= 8'h97;
         1779: data_out <= 8'h9e;
         1780: data_out <= 8'hbd;
         1781: data_out <= 8'h02;
         1782: data_out <= 8'hb5;
         1783: data_out <= 8'h35;
         1784: data_out <= 8'h81;
         1785: data_out <= 8'h0b;
         1786: data_out <= 8'h27;
         1787: data_out <= 8'h0b;
         1788: data_out <= 8'hc6;
         1789: data_out <= 8'h04;
         1790: data_out <= 8'h8c;
         1791: data_out <= 8'hc6;
         1792: data_out <= 8'h0e;
         1793: data_out <= 8'h7e;
         1794: data_out <= 8'h03;
         1795: data_out <= 8'h21;
         1796: data_out <= 8'h7e;
         1797: data_out <= 8'h0b;
         1798: data_out <= 8'h57;
         1799: data_out <= 8'h32;
         1800: data_out <= 8'h33;
         1801: data_out <= 8'hd7;
         1802: data_out <= 8'h8a;
         1803: data_out <= 8'h33;
         1804: data_out <= 8'hd7;
         1805: data_out <= 8'h8b;
         1806: data_out <= 8'h33;
         1807: data_out <= 8'hd7;
         1808: data_out <= 8'hc8;
         1809: data_out <= 8'h33;
         1810: data_out <= 8'hd7;
         1811: data_out <= 8'hc9;
         1812: data_out <= 8'h8d;
         1813: data_out <= 8'h03;
         1814: data_out <= 8'hdf;
         1815: data_out <= 8'hc8;
         1816: data_out <= 8'h39;
         1817: data_out <= 8'hc6;
         1818: data_out <= 8'h3a;
         1819: data_out <= 8'h86;
         1820: data_out <= 8'h5f;
         1821: data_out <= 8'hd7;
         1822: data_out <= 8'h58;
         1823: data_out <= 8'h5f;
         1824: data_out <= 8'hde;
         1825: data_out <= 8'hc8;
         1826: data_out <= 8'h17;
         1827: data_out <= 8'hd6;
         1828: data_out <= 8'h58;
         1829: data_out <= 8'h97;
         1830: data_out <= 8'h58;
         1831: data_out <= 8'ha6;
         1832: data_out <= 8'h00;
         1833: data_out <= 8'h27;
         1834: data_out <= 8'hed;
         1835: data_out <= 8'h11;
         1836: data_out <= 8'h27;
         1837: data_out <= 8'hea;
         1838: data_out <= 8'h08;
         1839: data_out <= 8'h81;
         1840: data_out <= 8'h22;
         1841: data_out <= 8'h27;
         1842: data_out <= 8'hef;
         1843: data_out <= 8'h20;
         1844: data_out <= 8'hf2;
         1845: data_out <= 8'hbd;
         1846: data_out <= 8'h0a;
         1847: data_out <= 8'h27;
         1848: data_out <= 8'hbd;
         1849: data_out <= 8'h00;
         1850: data_out <= 8'hc7;
         1851: data_out <= 8'h81;
         1852: data_out <= 8'h88;
         1853: data_out <= 8'h27;
         1854: data_out <= 8'h05;
         1855: data_out <= 8'hc6;
         1856: data_out <= 8'ha0;
         1857: data_out <= 8'hbd;
         1858: data_out <= 8'h0b;
         1859: data_out <= 8'h4d;
         1860: data_out <= 8'h96;
         1861: data_out <= 8'haf;
         1862: data_out <= 8'h26;
         1863: data_out <= 8'h05;
         1864: data_out <= 8'h8d;
         1865: data_out <= 8'hd2;
         1866: data_out <= 8'hdf;
         1867: data_out <= 8'hc8;
         1868: data_out <= 8'h39;
         1869: data_out <= 8'hbd;
         1870: data_out <= 8'h00;
         1871: data_out <= 8'hc7;
         1872: data_out <= 8'h25;
         1873: data_out <= 8'h85;
         1874: data_out <= 8'h7e;
         1875: data_out <= 8'h06;
         1876: data_out <= 8'h04;
         1877: data_out <= 8'hbd;
         1878: data_out <= 8'h11;
         1879: data_out <= 8'h6a;
         1880: data_out <= 8'h36;
         1881: data_out <= 8'h81;
         1882: data_out <= 8'h8c;
         1883: data_out <= 8'h27;
         1884: data_out <= 8'h04;
         1885: data_out <= 8'h81;
         1886: data_out <= 8'h88;
         1887: data_out <= 8'h26;
         1888: data_out <= 8'ha3;
         1889: data_out <= 8'h7a;
         1890: data_out <= 8'h00;
         1891: data_out <= 8'hb2;
         1892: data_out <= 8'h26;
         1893: data_out <= 8'h04;
         1894: data_out <= 8'h32;
         1895: data_out <= 8'h7e;
         1896: data_out <= 8'h06;
         1897: data_out <= 8'h06;
         1898: data_out <= 8'hbd;
         1899: data_out <= 8'h00;
         1900: data_out <= 8'hbf;
         1901: data_out <= 8'h8d;
         1902: data_out <= 8'h06;
         1903: data_out <= 8'h81;
         1904: data_out <= 8'h2c;
         1905: data_out <= 8'h27;
         1906: data_out <= 8'hee;
         1907: data_out <= 8'h31;
         1908: data_out <= 8'h39;
         1909: data_out <= 8'hce;
         1910: data_out <= 8'h00;
         1911: data_out <= 8'h00;
         1912: data_out <= 8'hdf;
         1913: data_out <= 8'h8e;
         1914: data_out <= 8'h24;
         1915: data_out <= 8'hf8;
         1916: data_out <= 8'h80;
         1917: data_out <= 8'h30;
         1918: data_out <= 8'h97;
         1919: data_out <= 8'h58;
         1920: data_out <= 8'h96;
         1921: data_out <= 8'h8e;
         1922: data_out <= 8'hd6;
         1923: data_out <= 8'h8f;
         1924: data_out <= 8'h81;
         1925: data_out <= 8'h18;
         1926: data_out <= 8'h22;
         1927: data_out <= 8'hd7;
         1928: data_out <= 8'h58;
         1929: data_out <= 8'h49;
         1930: data_out <= 8'h58;
         1931: data_out <= 8'h49;
         1932: data_out <= 8'hdb;
         1933: data_out <= 8'h8f;
         1934: data_out <= 8'h99;
         1935: data_out <= 8'h8e;
         1936: data_out <= 8'h58;
         1937: data_out <= 8'h49;
         1938: data_out <= 8'hdb;
         1939: data_out <= 8'h58;
         1940: data_out <= 8'h89;
         1941: data_out <= 8'h00;
         1942: data_out <= 8'h97;
         1943: data_out <= 8'h8e;
         1944: data_out <= 8'hd7;
         1945: data_out <= 8'h8f;
         1946: data_out <= 8'hbd;
         1947: data_out <= 8'h00;
         1948: data_out <= 8'hbf;
         1949: data_out <= 8'h20;
         1950: data_out <= 8'hdb;
         1951: data_out <= 8'hbd;
         1952: data_out <= 8'h0c;
         1953: data_out <= 8'h37;
         1954: data_out <= 8'hdf;
         1955: data_out <= 8'h9e;
         1956: data_out <= 8'hc6;
         1957: data_out <= 8'hab;
         1958: data_out <= 8'hbd;
         1959: data_out <= 8'h0b;
         1960: data_out <= 8'h4d;
         1961: data_out <= 8'h96;
         1962: data_out <= 8'h5c;
         1963: data_out <= 8'h36;
         1964: data_out <= 8'hbd;
         1965: data_out <= 8'h0a;
         1966: data_out <= 8'h27;
         1967: data_out <= 8'h32;
         1968: data_out <= 8'h46;
         1969: data_out <= 8'hbd;
         1970: data_out <= 8'h0a;
         1971: data_out <= 8'h1d;
         1972: data_out <= 8'h27;
         1973: data_out <= 8'h49;
         1974: data_out <= 8'hde;
         1975: data_out <= 8'hb1;
         1976: data_out <= 8'h96;
         1977: data_out <= 8'h82;
         1978: data_out <= 8'ha1;
         1979: data_out <= 8'h02;
         1980: data_out <= 8'h22;
         1981: data_out <= 8'h23;
         1982: data_out <= 8'h25;
         1983: data_out <= 8'h06;
         1984: data_out <= 8'hd6;
         1985: data_out <= 8'h83;
         1986: data_out <= 8'he1;
         1987: data_out <= 8'h03;
         1988: data_out <= 8'h24;
         1989: data_out <= 8'h1b;
         1990: data_out <= 8'h96;
         1991: data_out <= 8'h7c;
         1992: data_out <= 8'h91;
         1993: data_out <= 8'hb1;
         1994: data_out <= 8'h22;
         1995: data_out <= 8'h15;
         1996: data_out <= 8'h25;
         1997: data_out <= 8'h06;
         1998: data_out <= 8'hd6;
         1999: data_out <= 8'h7c;
         2000: data_out <= 8'hd1;
         2001: data_out <= 8'hb2;
         2002: data_out <= 8'h22;
         2003: data_out <= 8'h0d;
         2004: data_out <= 8'he6;
         2005: data_out <= 8'h00;
         2006: data_out <= 8'hbd;
         2007: data_out <= 8'h0f;
         2008: data_out <= 8'h2d;
         2009: data_out <= 8'hde;
         2010: data_out <= 8'had;
         2011: data_out <= 8'hbd;
         2012: data_out <= 8'h10;
         2013: data_out <= 8'h8b;
         2014: data_out <= 8'hce;
         2015: data_out <= 8'h00;
         2016: data_out <= 8'haf;
         2017: data_out <= 8'hdf;
         2018: data_out <= 8'had;
         2019: data_out <= 8'hbd;
         2020: data_out <= 8'h10;
         2021: data_out <= 8'hc7;
         2022: data_out <= 8'h07;
         2023: data_out <= 8'h36;
         2024: data_out <= 8'h9f;
         2025: data_out <= 8'h78;
         2026: data_out <= 8'h0f;
         2027: data_out <= 8'hde;
         2028: data_out <= 8'had;
         2029: data_out <= 8'h35;
         2030: data_out <= 8'hde;
         2031: data_out <= 8'h9e;
         2032: data_out <= 8'h32;
         2033: data_out <= 8'ha7;
         2034: data_out <= 8'h00;
         2035: data_out <= 8'h32;
         2036: data_out <= 8'h32;
         2037: data_out <= 8'ha7;
         2038: data_out <= 8'h02;
         2039: data_out <= 8'h32;
         2040: data_out <= 8'ha7;
         2041: data_out <= 8'h03;
         2042: data_out <= 8'h9e;
         2043: data_out <= 8'h78;
         2044: data_out <= 8'h32;
         2045: data_out <= 8'h06;
         2046: data_out <= 8'h39;
         2047: data_out <= 8'h7e;
         2048: data_out <= 8'h15;
         2049: data_out <= 8'ha8;
         2050: data_out <= 8'hbd;
         2051: data_out <= 8'h08;
         2052: data_out <= 8'h8a;
         2053: data_out <= 8'hbd;
         2054: data_out <= 8'h00;
         2055: data_out <= 8'hc7;
         2056: data_out <= 8'h27;
         2057: data_out <= 8'h38;
         2058: data_out <= 8'h27;
         2059: data_out <= 8'h4e;
         2060: data_out <= 8'h81;
         2061: data_out <= 8'h9c;
         2062: data_out <= 8'h27;
         2063: data_out <= 8'h5c;
         2064: data_out <= 8'h81;
         2065: data_out <= 8'h9f;
         2066: data_out <= 8'h27;
         2067: data_out <= 8'h58;
         2068: data_out <= 8'h81;
         2069: data_out <= 8'h2c;
         2070: data_out <= 8'h27;
         2071: data_out <= 8'h43;
         2072: data_out <= 8'h81;
         2073: data_out <= 8'h3b;
         2074: data_out <= 8'h27;
         2075: data_out <= 8'h66;
         2076: data_out <= 8'hbd;
         2077: data_out <= 8'h0a;
         2078: data_out <= 8'h27;
         2079: data_out <= 8'hde;
         2080: data_out <= 8'hb1;
         2081: data_out <= 8'h96;
         2082: data_out <= 8'h5c;
         2083: data_out <= 8'h26;
         2084: data_out <= 8'hdd;
         2085: data_out <= 8'hbd;
         2086: data_out <= 8'h17;
         2087: data_out <= 8'h45;
         2088: data_out <= 8'hbd;
         2089: data_out <= 8'h0f;
         2090: data_out <= 8'h36;
         2091: data_out <= 8'hde;
         2092: data_out <= 8'hb1;
         2093: data_out <= 8'h96;
         2094: data_out <= 8'h0b;
         2095: data_out <= 8'hab;
         2096: data_out <= 8'h00;
         2097: data_out <= 8'h91;
         2098: data_out <= 8'h0c;
         2099: data_out <= 8'h23;
         2100: data_out <= 8'h02;
         2101: data_out <= 8'h8d;
         2102: data_out <= 8'h0b;
         2103: data_out <= 8'h8d;
         2104: data_out <= 8'h51;
         2105: data_out <= 8'h8d;
         2106: data_out <= 8'h63;
         2107: data_out <= 8'h20;
         2108: data_out <= 8'hc8;
         2109: data_out <= 8'h6f;
         2110: data_out <= 8'h00;
         2111: data_out <= 8'hce;
         2112: data_out <= 8'h00;
         2113: data_out <= 8'h0f;
         2114: data_out <= 8'h86;
         2115: data_out <= 8'h0d;
         2116: data_out <= 8'h97;
         2117: data_out <= 8'h0b;
         2118: data_out <= 8'h8d;
         2119: data_out <= 8'h5b;
         2120: data_out <= 8'h86;
         2121: data_out <= 8'h0a;
         2122: data_out <= 8'h8d;
         2123: data_out <= 8'h57;
         2124: data_out <= 8'h37;
         2125: data_out <= 8'hd6;
         2126: data_out <= 8'h0a;
         2127: data_out <= 8'h27;
         2128: data_out <= 8'h06;
         2129: data_out <= 8'h4f;
         2130: data_out <= 8'h8d;
         2131: data_out <= 8'h4f;
         2132: data_out <= 8'h5a;
         2133: data_out <= 8'h26;
         2134: data_out <= 8'hfb;
         2135: data_out <= 8'hd7;
         2136: data_out <= 8'h0b;
         2137: data_out <= 8'h33;
         2138: data_out <= 8'h39;
         2139: data_out <= 8'hd6;
         2140: data_out <= 8'h0b;
         2141: data_out <= 8'hd1;
         2142: data_out <= 8'h0d;
         2143: data_out <= 8'h25;
         2144: data_out <= 8'h04;
         2145: data_out <= 8'h8d;
         2146: data_out <= 8'hdf;
         2147: data_out <= 8'h20;
         2148: data_out <= 8'h1d;
         2149: data_out <= 8'hc0;
         2150: data_out <= 8'h0e;
         2151: data_out <= 8'h24;
         2152: data_out <= 8'hfc;
         2153: data_out <= 8'h50;
         2154: data_out <= 8'h20;
         2155: data_out <= 8'h11;
         2156: data_out <= 8'h36;
         2157: data_out <= 8'hbd;
         2158: data_out <= 8'h11;
         2159: data_out <= 8'h67;
         2160: data_out <= 8'h81;
         2161: data_out <= 8'h29;
         2162: data_out <= 8'h26;
         2163: data_out <= 8'h67;
         2164: data_out <= 8'h32;
         2165: data_out <= 8'h81;
         2166: data_out <= 8'h9f;
         2167: data_out <= 8'h27;
         2168: data_out <= 8'h04;
         2169: data_out <= 8'hd0;
         2170: data_out <= 8'h0b;
         2171: data_out <= 8'h23;
         2172: data_out <= 8'h05;
         2173: data_out <= 8'h8d;
         2174: data_out <= 8'h1f;
         2175: data_out <= 8'h5a;
         2176: data_out <= 8'h26;
         2177: data_out <= 8'hfb;
         2178: data_out <= 8'hbd;
         2179: data_out <= 8'h00;
         2180: data_out <= 8'hbf;
         2181: data_out <= 8'h20;
         2182: data_out <= 8'h83;
         2183: data_out <= 8'hbd;
         2184: data_out <= 8'h0f;
         2185: data_out <= 8'h37;
         2186: data_out <= 8'hbd;
         2187: data_out <= 8'h10;
         2188: data_out <= 8'ha9;
         2189: data_out <= 8'h5c;
         2190: data_out <= 8'h5a;
         2191: data_out <= 8'h27;
         2192: data_out <= 8'hc9;
         2193: data_out <= 8'ha6;
         2194: data_out <= 8'h00;
         2195: data_out <= 8'h8d;
         2196: data_out <= 8'h0e;
         2197: data_out <= 8'h08;
         2198: data_out <= 8'h81;
         2199: data_out <= 8'h0d;
         2200: data_out <= 8'h26;
         2201: data_out <= 8'hf4;
         2202: data_out <= 8'h8d;
         2203: data_out <= 8'hb0;
         2204: data_out <= 8'h20;
         2205: data_out <= 8'hf0;
         2206: data_out <= 8'h86;
         2207: data_out <= 8'h20;
         2208: data_out <= 8'h8c;
         2209: data_out <= 8'h86;
         2210: data_out <= 8'h3f;
         2211: data_out <= 8'h7d;
         2212: data_out <= 8'h01;
         2213: data_out <= 8'h11;
         2214: data_out <= 8'h26;
         2215: data_out <= 8'h17;
         2216: data_out <= 8'h36;
         2217: data_out <= 8'h81;
         2218: data_out <= 8'h20;
         2219: data_out <= 8'h25;
         2220: data_out <= 8'h0b;
         2221: data_out <= 8'h96;
         2222: data_out <= 8'h0b;
         2223: data_out <= 8'h91;
         2224: data_out <= 8'h0c;
         2225: data_out <= 8'h26;
         2226: data_out <= 8'h02;
         2227: data_out <= 8'h8d;
         2228: data_out <= 8'h8d;
         2229: data_out <= 8'h4c;
         2230: data_out <= 8'h97;
         2231: data_out <= 8'h0b;
         2232: data_out <= 8'h32;
         2233: data_out <= 8'h37;
         2234: data_out <= 8'h16;
         2235: data_out <= 8'hbd;
         2236: data_out <= 8'hff;
         2237: data_out <= 8'h81;
         2238: data_out <= 8'h33;
         2239: data_out <= 8'h39;
         2240: data_out <= 8'h3f;
         2241: data_out <= 8'h52;
         2242: data_out <= 8'h45;
         2243: data_out <= 8'h44;
         2244: data_out <= 8'h4f;
         2245: data_out <= 8'h20;
         2246: data_out <= 8'h46;
         2247: data_out <= 8'h52;
         2248: data_out <= 8'h4f;
         2249: data_out <= 8'h4d;
         2250: data_out <= 8'h20;
         2251: data_out <= 8'h53;
         2252: data_out <= 8'h54;
         2253: data_out <= 8'h41;
         2254: data_out <= 8'h52;
         2255: data_out <= 8'hd4;
         2256: data_out <= 8'h0d;
         2257: data_out <= 8'h0a;
         2258: data_out <= 8'h00;
         2259: data_out <= 8'h96;
         2260: data_out <= 8'h5f;
         2261: data_out <= 8'h27;
         2262: data_out <= 8'h07;
         2263: data_out <= 8'hde;
         2264: data_out <= 8'h94;
         2265: data_out <= 8'hdf;
         2266: data_out <= 8'h8a;
         2267: data_out <= 8'h7e;
         2268: data_out <= 8'h0b;
         2269: data_out <= 8'h57;
         2270: data_out <= 8'hce;
         2271: data_out <= 8'h08;
         2272: data_out <= 8'hbf;
         2273: data_out <= 8'h8d;
         2274: data_out <= 8'ha4;
         2275: data_out <= 8'hde;
         2276: data_out <= 8'h92;
         2277: data_out <= 8'hdf;
         2278: data_out <= 8'hc8;
         2279: data_out <= 8'h39;
         2280: data_out <= 8'h7f;
         2281: data_out <= 8'h01;
         2282: data_out <= 8'h11;
         2283: data_out <= 8'h81;
         2284: data_out <= 8'h22;
         2285: data_out <= 8'h26;
         2286: data_out <= 8'h0a;
         2287: data_out <= 8'hbd;
         2288: data_out <= 8'h0b;
         2289: data_out <= 8'h18;
         2290: data_out <= 8'hc6;
         2291: data_out <= 8'h3b;
         2292: data_out <= 8'hbd;
         2293: data_out <= 8'h0b;
         2294: data_out <= 8'h4d;
         2295: data_out <= 8'h8d;
         2296: data_out <= 8'h91;
         2297: data_out <= 8'hbd;
         2298: data_out <= 8'h0e;
         2299: data_out <= 8'h71;
         2300: data_out <= 8'h8d;
         2301: data_out <= 8'h09;
         2302: data_out <= 8'h96;
         2303: data_out <= 8'h10;
         2304: data_out <= 8'h26;
         2305: data_out <= 8'h0f;
         2306: data_out <= 8'h0c;
         2307: data_out <= 8'h07;
         2308: data_out <= 8'h7e;
         2309: data_out <= 8'h06;
         2310: data_out <= 8'h43;
         2311: data_out <= 8'h8d;
         2312: data_out <= 8'h98;
         2313: data_out <= 8'h8d;
         2314: data_out <= 8'h93;
         2315: data_out <= 8'h7e;
         2316: data_out <= 8'h03;
         2317: data_out <= 8'hfa;
         2318: data_out <= 8'hde;
         2319: data_out <= 8'h96;
         2320: data_out <= 8'h86;
         2321: data_out <= 8'h4f;
         2322: data_out <= 8'h97;
         2323: data_out <= 8'h5f;
         2324: data_out <= 8'hdf;
         2325: data_out <= 8'h98;
         2326: data_out <= 8'hbd;
         2327: data_out <= 8'h0c;
         2328: data_out <= 8'h37;
         2329: data_out <= 8'hdf;
         2330: data_out <= 8'h9e;
         2331: data_out <= 8'hde;
         2332: data_out <= 8'hc8;
         2333: data_out <= 8'hdf;
         2334: data_out <= 8'h8e;
         2335: data_out <= 8'hde;
         2336: data_out <= 8'h98;
         2337: data_out <= 8'ha6;
         2338: data_out <= 8'h00;
         2339: data_out <= 8'h26;
         2340: data_out <= 8'h09;
         2341: data_out <= 8'h96;
         2342: data_out <= 8'h5f;
         2343: data_out <= 8'h26;
         2344: data_out <= 8'h4e;
         2345: data_out <= 8'hbd;
         2346: data_out <= 8'h08;
         2347: data_out <= 8'ha1;
         2348: data_out <= 8'h8d;
         2349: data_out <= 8'hd9;
         2350: data_out <= 8'hdf;
         2351: data_out <= 8'hc8;
         2352: data_out <= 8'hbd;
         2353: data_out <= 8'h00;
         2354: data_out <= 8'hbf;
         2355: data_out <= 8'hd6;
         2356: data_out <= 8'h5c;
         2357: data_out <= 8'h27;
         2358: data_out <= 8'h1c;
         2359: data_out <= 8'hde;
         2360: data_out <= 8'hc8;
         2361: data_out <= 8'h97;
         2362: data_out <= 8'h58;
         2363: data_out <= 8'h81;
         2364: data_out <= 8'h22;
         2365: data_out <= 8'h27;
         2366: data_out <= 8'h07;
         2367: data_out <= 8'h09;
         2368: data_out <= 8'h86;
         2369: data_out <= 8'h3a;
         2370: data_out <= 8'h97;
         2371: data_out <= 8'h58;
         2372: data_out <= 8'h86;
         2373: data_out <= 8'h2c;
         2374: data_out <= 8'h97;
         2375: data_out <= 8'h59;
         2376: data_out <= 8'hbd;
         2377: data_out <= 8'h0f;
         2378: data_out <= 8'h3d;
         2379: data_out <= 8'hbd;
         2380: data_out <= 8'h11;
         2381: data_out <= 8'h9b;
         2382: data_out <= 8'hbd;
         2383: data_out <= 8'h07;
         2384: data_out <= 8'hb6;
         2385: data_out <= 8'h20;
         2386: data_out <= 8'h06;
         2387: data_out <= 8'hbd;
         2388: data_out <= 8'h16;
         2389: data_out <= 8'h7c;
         2390: data_out <= 8'hbd;
         2391: data_out <= 8'h15;
         2392: data_out <= 8'ha8;
         2393: data_out <= 8'hbd;
         2394: data_out <= 8'h00;
         2395: data_out <= 8'hc7;
         2396: data_out <= 8'h27;
         2397: data_out <= 8'h07;
         2398: data_out <= 8'h81;
         2399: data_out <= 8'h2c;
         2400: data_out <= 8'h27;
         2401: data_out <= 8'h03;
         2402: data_out <= 8'h7e;
         2403: data_out <= 8'h08;
         2404: data_out <= 8'hd3;
         2405: data_out <= 8'hde;
         2406: data_out <= 8'hc8;
         2407: data_out <= 8'hdf;
         2408: data_out <= 8'h98;
         2409: data_out <= 8'hde;
         2410: data_out <= 8'h8e;
         2411: data_out <= 8'hdf;
         2412: data_out <= 8'hc8;
         2413: data_out <= 8'hbd;
         2414: data_out <= 8'h00;
         2415: data_out <= 8'hc7;
         2416: data_out <= 8'h27;
         2417: data_out <= 8'h2a;
         2418: data_out <= 8'hbd;
         2419: data_out <= 8'h0b;
         2420: data_out <= 8'h4b;
         2421: data_out <= 8'h20;
         2422: data_out <= 8'h9f;
         2423: data_out <= 8'hdf;
         2424: data_out <= 8'hc8;
         2425: data_out <= 8'hbd;
         2426: data_out <= 8'h07;
         2427: data_out <= 8'h19;
         2428: data_out <= 8'h4d;
         2429: data_out <= 8'h26;
         2430: data_out <= 8'h14;
         2431: data_out <= 8'ha6;
         2432: data_out <= 8'h01;
         2433: data_out <= 8'hc6;
         2434: data_out <= 8'h06;
         2435: data_out <= 8'haa;
         2436: data_out <= 8'h02;
         2437: data_out <= 8'h27;
         2438: data_out <= 8'h4d;
         2439: data_out <= 8'ha6;
         2440: data_out <= 8'h03;
         2441: data_out <= 8'h97;
         2442: data_out <= 8'h94;
         2443: data_out <= 8'ha6;
         2444: data_out <= 8'h04;
         2445: data_out <= 8'h97;
         2446: data_out <= 8'h95;
         2447: data_out <= 8'h08;
         2448: data_out <= 8'h08;
         2449: data_out <= 8'h08;
         2450: data_out <= 8'h08;
         2451: data_out <= 8'h08;
         2452: data_out <= 8'ha6;
         2453: data_out <= 8'h00;
         2454: data_out <= 8'h81;
         2455: data_out <= 8'h83;
         2456: data_out <= 8'h26;
         2457: data_out <= 8'hdd;
         2458: data_out <= 8'h20;
         2459: data_out <= 8'h92;
         2460: data_out <= 8'hde;
         2461: data_out <= 8'h98;
         2462: data_out <= 8'hd6;
         2463: data_out <= 8'h5f;
         2464: data_out <= 8'h27;
         2465: data_out <= 8'h03;
         2466: data_out <= 8'h7e;
         2467: data_out <= 8'h06;
         2468: data_out <= 8'h23;
         2469: data_out <= 8'ha6;
         2470: data_out <= 8'h00;
         2471: data_out <= 8'h27;
         2472: data_out <= 8'h06;
         2473: data_out <= 8'hce;
         2474: data_out <= 8'h09;
         2475: data_out <= 8'haf;
         2476: data_out <= 8'h7e;
         2477: data_out <= 8'h08;
         2478: data_out <= 8'h87;
         2479: data_out <= 8'h39;
         2480: data_out <= 8'h3f;
         2481: data_out <= 8'h45;
         2482: data_out <= 8'h58;
         2483: data_out <= 8'h54;
         2484: data_out <= 8'h52;
         2485: data_out <= 8'h41;
         2486: data_out <= 8'h20;
         2487: data_out <= 8'h49;
         2488: data_out <= 8'h47;
         2489: data_out <= 8'h4e;
         2490: data_out <= 8'h4f;
         2491: data_out <= 8'h52;
         2492: data_out <= 8'h45;
         2493: data_out <= 8'hc4;
         2494: data_out <= 8'h0d;
         2495: data_out <= 8'h0a;
         2496: data_out <= 8'h00;
         2497: data_out <= 8'h26;
         2498: data_out <= 8'h05;
         2499: data_out <= 8'hce;
         2500: data_out <= 8'h00;
         2501: data_out <= 8'h00;
         2502: data_out <= 8'h20;
         2503: data_out <= 8'h03;
         2504: data_out <= 8'hbd;
         2505: data_out <= 8'h0c;
         2506: data_out <= 8'h37;
         2507: data_out <= 8'hdf;
         2508: data_out <= 8'h9e;
         2509: data_out <= 8'hbd;
         2510: data_out <= 8'h02;
         2511: data_out <= 8'hb5;
         2512: data_out <= 8'h27;
         2513: data_out <= 8'h04;
         2514: data_out <= 8'hc6;
         2515: data_out <= 8'h00;
         2516: data_out <= 8'h20;
         2517: data_out <= 8'h4e;
         2518: data_out <= 8'h35;
         2519: data_out <= 8'h08;
         2520: data_out <= 8'h08;
         2521: data_out <= 8'h08;
         2522: data_out <= 8'hdf;
         2523: data_out <= 8'h71;
         2524: data_out <= 8'hbd;
         2525: data_out <= 8'h15;
         2526: data_out <= 8'h8e;
         2527: data_out <= 8'h30;
         2528: data_out <= 8'ha6;
         2529: data_out <= 8'h07;
         2530: data_out <= 8'h97;
         2531: data_out <= 8'hb3;
         2532: data_out <= 8'hde;
         2533: data_out <= 8'h9e;
         2534: data_out <= 8'hbd;
         2535: data_out <= 8'h13;
         2536: data_out <= 8'h1a;
         2537: data_out <= 8'hbd;
         2538: data_out <= 8'h15;
         2539: data_out <= 8'ha8;
         2540: data_out <= 8'hde;
         2541: data_out <= 8'h71;
         2542: data_out <= 8'h08;
         2543: data_out <= 8'h08;
         2544: data_out <= 8'h08;
         2545: data_out <= 8'h08;
         2546: data_out <= 8'h08;
         2547: data_out <= 8'hbd;
         2548: data_out <= 8'h16;
         2549: data_out <= 8'h04;
         2550: data_out <= 8'h30;
         2551: data_out <= 8'he0;
         2552: data_out <= 8'h07;
         2553: data_out <= 8'h27;
         2554: data_out <= 8'h0c;
         2555: data_out <= 8'hee;
         2556: data_out <= 8'h0c;
         2557: data_out <= 8'hdf;
         2558: data_out <= 8'h8a;
         2559: data_out <= 8'h30;
         2560: data_out <= 8'hee;
         2561: data_out <= 8'h0e;
         2562: data_out <= 8'hdf;
         2563: data_out <= 8'hc8;
         2564: data_out <= 8'h7e;
         2565: data_out <= 8'h05;
         2566: data_out <= 8'hd6;
         2567: data_out <= 8'hc6;
         2568: data_out <= 8'h10;
         2569: data_out <= 8'hbd;
         2570: data_out <= 8'h03;
         2571: data_out <= 8'h11;
         2572: data_out <= 8'h35;
         2573: data_out <= 8'hbd;
         2574: data_out <= 8'h00;
         2575: data_out <= 8'hc7;
         2576: data_out <= 8'h81;
         2577: data_out <= 8'h2c;
         2578: data_out <= 8'h26;
         2579: data_out <= 8'hf0;
         2580: data_out <= 8'hbd;
         2581: data_out <= 8'h00;
         2582: data_out <= 8'hbf;
         2583: data_out <= 8'h8d;
         2584: data_out <= 8'haf;
         2585: data_out <= 8'h8d;
         2586: data_out <= 8'h0c;
         2587: data_out <= 8'h6d;
         2588: data_out <= 8'h0d;
         2589: data_out <= 8'h76;
         2590: data_out <= 8'h00;
         2591: data_out <= 8'h5c;
         2592: data_out <= 8'h28;
         2593: data_out <= 8'h8d;
         2594: data_out <= 8'hc6;
         2595: data_out <= 8'h18;
         2596: data_out <= 8'h7e;
         2597: data_out <= 8'h03;
         2598: data_out <= 8'h21;
         2599: data_out <= 8'hde;
         2600: data_out <= 8'hc8;
         2601: data_out <= 8'h09;
         2602: data_out <= 8'hdf;
         2603: data_out <= 8'hc8;
         2604: data_out <= 8'h4f;
         2605: data_out <= 8'hc6;
         2606: data_out <= 8'h37;
         2607: data_out <= 8'h36;
         2608: data_out <= 8'hc6;
         2609: data_out <= 8'h01;
         2610: data_out <= 8'hbd;
         2611: data_out <= 8'h02;
         2612: data_out <= 8'hf8;
         2613: data_out <= 8'hbd;
         2614: data_out <= 8'h0a;
         2615: data_out <= 8'hf9;
         2616: data_out <= 8'h7f;
         2617: data_out <= 8'h00;
         2618: data_out <= 8'ha2;
         2619: data_out <= 8'hbd;
         2620: data_out <= 8'h00;
         2621: data_out <= 8'hc7;
         2622: data_out <= 8'h80;
         2623: data_out <= 8'haa;
         2624: data_out <= 8'h25;
         2625: data_out <= 8'h14;
         2626: data_out <= 8'h81;
         2627: data_out <= 8'h03;
         2628: data_out <= 8'h24;
         2629: data_out <= 8'h10;
         2630: data_out <= 8'h81;
         2631: data_out <= 8'h01;
         2632: data_out <= 8'h49;
         2633: data_out <= 8'h98;
         2634: data_out <= 8'ha2;
         2635: data_out <= 8'h91;
         2636: data_out <= 8'ha2;
         2637: data_out <= 8'h25;
         2638: data_out <= 8'h5d;
         2639: data_out <= 8'h97;
         2640: data_out <= 8'ha2;
         2641: data_out <= 8'hbd;
         2642: data_out <= 8'h00;
         2643: data_out <= 8'hbf;
         2644: data_out <= 8'h20;
         2645: data_out <= 8'he8;
         2646: data_out <= 8'hd6;
         2647: data_out <= 8'ha2;
         2648: data_out <= 8'h26;
         2649: data_out <= 8'h2d;
         2650: data_out <= 8'h24;
         2651: data_out <= 8'h6b;
         2652: data_out <= 8'h8b;
         2653: data_out <= 8'h07;
         2654: data_out <= 8'h24;
         2655: data_out <= 8'h67;
         2656: data_out <= 8'h99;
         2657: data_out <= 8'h5c;
         2658: data_out <= 8'h26;
         2659: data_out <= 8'h03;
         2660: data_out <= 8'h7e;
         2661: data_out <= 8'h10;
         2662: data_out <= 8'h51;
         2663: data_out <= 8'h89;
         2664: data_out <= 8'hff;
         2665: data_out <= 8'h16;
         2666: data_out <= 8'h48;
         2667: data_out <= 8'h1b;
         2668: data_out <= 8'h16;
         2669: data_out <= 8'hce;
         2670: data_out <= 8'h01;
         2671: data_out <= 8'h47;
         2672: data_out <= 8'hbd;
         2673: data_out <= 8'h03;
         2674: data_out <= 8'h11;
         2675: data_out <= 8'h32;
         2676: data_out <= 8'ha1;
         2677: data_out <= 8'h00;
         2678: data_out <= 8'h24;
         2679: data_out <= 8'h56;
         2680: data_out <= 8'h8d;
         2681: data_out <= 8'ha1;
         2682: data_out <= 8'h36;
         2683: data_out <= 8'h8d;
         2684: data_out <= 8'h23;
         2685: data_out <= 8'hde;
         2686: data_out <= 8'ha0;
         2687: data_out <= 8'h32;
         2688: data_out <= 8'h26;
         2689: data_out <= 8'h18;
         2690: data_out <= 8'h4d;
         2691: data_out <= 8'h27;
         2692: data_out <= 8'h71;
         2693: data_out <= 8'h20;
         2694: data_out <= 8'h50;
         2695: data_out <= 8'h78;
         2696: data_out <= 8'h00;
         2697: data_out <= 8'h5c;
         2698: data_out <= 8'h59;
         2699: data_out <= 8'hde;
         2700: data_out <= 8'hc8;
         2701: data_out <= 8'h09;
         2702: data_out <= 8'hdf;
         2703: data_out <= 8'hc8;
         2704: data_out <= 8'hce;
         2705: data_out <= 8'h0a;
         2706: data_out <= 8'h97;
         2707: data_out <= 8'hd7;
         2708: data_out <= 8'ha2;
         2709: data_out <= 8'h20;
         2710: data_out <= 8'hdc;
         2711: data_out <= 8'h64;
         2712: data_out <= 8'h0b;
         2713: data_out <= 8'hca;
         2714: data_out <= 8'ha1;
         2715: data_out <= 8'h00;
         2716: data_out <= 8'h24;
         2717: data_out <= 8'h39;
         2718: data_out <= 8'h20;
         2719: data_out <= 8'hda;
         2720: data_out <= 8'ha6;
         2721: data_out <= 8'h02;
         2722: data_out <= 8'h36;
         2723: data_out <= 8'ha6;
         2724: data_out <= 8'h01;
         2725: data_out <= 8'h36;
         2726: data_out <= 8'h8d;
         2727: data_out <= 8'h07;
         2728: data_out <= 8'hd6;
         2729: data_out <= 8'ha2;
         2730: data_out <= 8'h20;
         2731: data_out <= 8'h82;
         2732: data_out <= 8'h7e;
         2733: data_out <= 8'h0b;
         2734: data_out <= 8'h57;
         2735: data_out <= 8'hd6;
         2736: data_out <= 8'hb3;
         2737: data_out <= 8'ha6;
         2738: data_out <= 8'h00;
         2739: data_out <= 8'h30;
         2740: data_out <= 8'hee;
         2741: data_out <= 8'h00;
         2742: data_out <= 8'h31;
         2743: data_out <= 8'h31;
         2744: data_out <= 8'h37;
         2745: data_out <= 8'hd6;
         2746: data_out <= 8'hb2;
         2747: data_out <= 8'h37;
         2748: data_out <= 8'hd6;
         2749: data_out <= 8'hb1;
         2750: data_out <= 8'h37;
         2751: data_out <= 8'hd6;
         2752: data_out <= 8'hb0;
         2753: data_out <= 8'h37;
         2754: data_out <= 8'hd6;
         2755: data_out <= 8'haf;
         2756: data_out <= 8'h37;
         2757: data_out <= 8'h6e;
         2758: data_out <= 8'h00;
         2759: data_out <= 8'hce;
         2760: data_out <= 8'h00;
         2761: data_out <= 8'h00;
         2762: data_out <= 8'h32;
         2763: data_out <= 8'h4d;
         2764: data_out <= 8'h27;
         2765: data_out <= 8'h28;
         2766: data_out <= 8'h81;
         2767: data_out <= 8'h64;
         2768: data_out <= 8'h27;
         2769: data_out <= 8'h03;
         2770: data_out <= 8'hbd;
         2771: data_out <= 8'h0a;
         2772: data_out <= 8'h1b;
         2773: data_out <= 8'hdf;
         2774: data_out <= 8'ha0;
         2775: data_out <= 8'h33;
         2776: data_out <= 8'h81;
         2777: data_out <= 8'h5a;
         2778: data_out <= 8'h27;
         2779: data_out <= 8'h1c;
         2780: data_out <= 8'h81;
         2781: data_out <= 8'h7d;
         2782: data_out <= 8'h27;
         2783: data_out <= 8'h18;
         2784: data_out <= 8'h54;
         2785: data_out <= 8'hd7;
         2786: data_out <= 8'h60;
         2787: data_out <= 8'h32;
         2788: data_out <= 8'h97;
         2789: data_out <= 8'hb6;
         2790: data_out <= 8'h33;
         2791: data_out <= 8'hd7;
         2792: data_out <= 8'hb7;
         2793: data_out <= 8'h33;
         2794: data_out <= 8'hd7;
         2795: data_out <= 8'hb8;
         2796: data_out <= 8'h33;
         2797: data_out <= 8'hd7;
         2798: data_out <= 8'hb9;
         2799: data_out <= 8'h33;
         2800: data_out <= 8'hd7;
         2801: data_out <= 8'hba;
         2802: data_out <= 8'hd8;
         2803: data_out <= 8'hb3;
         2804: data_out <= 8'hd7;
         2805: data_out <= 8'hbb;
         2806: data_out <= 8'hd6;
         2807: data_out <= 8'haf;
         2808: data_out <= 8'h39;
         2809: data_out <= 8'h7f;
         2810: data_out <= 8'h00;
         2811: data_out <= 8'h5c;
         2812: data_out <= 8'h8d;
         2813: data_out <= 8'h56;
         2814: data_out <= 8'h24;
         2815: data_out <= 8'h03;
         2816: data_out <= 8'h7e;
         2817: data_out <= 8'h16;
         2818: data_out <= 8'h7c;
         2819: data_out <= 8'hbd;
         2820: data_out <= 8'h0c;
         2821: data_out <= 8'h9b;
         2822: data_out <= 8'h24;
         2823: data_out <= 8'h5c;
         2824: data_out <= 8'h81;
         2825: data_out <= 8'h2e;
         2826: data_out <= 8'h27;
         2827: data_out <= 8'hf4;
         2828: data_out <= 8'h81;
         2829: data_out <= 8'ha4;
         2830: data_out <= 8'h27;
         2831: data_out <= 8'h4c;
         2832: data_out <= 8'h81;
         2833: data_out <= 8'ha3;
         2834: data_out <= 8'h27;
         2835: data_out <= 8'he8;
         2836: data_out <= 8'h81;
         2837: data_out <= 8'h22;
         2838: data_out <= 8'h26;
         2839: data_out <= 8'h08;
         2840: data_out <= 8'hde;
         2841: data_out <= 8'hc8;
         2842: data_out <= 8'hbd;
         2843: data_out <= 8'h0f;
         2844: data_out <= 8'h37;
         2845: data_out <= 8'h7e;
         2846: data_out <= 8'h11;
         2847: data_out <= 8'h9b;
         2848: data_out <= 8'h81;
         2849: data_out <= 8'ha1;
         2850: data_out <= 8'h26;
         2851: data_out <= 8'h11;
         2852: data_out <= 8'h86;
         2853: data_out <= 8'h5a;
         2854: data_out <= 8'hbd;
         2855: data_out <= 8'h0a;
         2856: data_out <= 8'h2e;
         2857: data_out <= 8'hbd;
         2858: data_out <= 8'h0c;
         2859: data_out <= 8'hf1;
         2860: data_out <= 8'h96;
         2861: data_out <= 8'hb1;
         2862: data_out <= 8'hd6;
         2863: data_out <= 8'hb2;
         2864: data_out <= 8'h43;
         2865: data_out <= 8'h53;
         2866: data_out <= 8'h7e;
         2867: data_out <= 8'h0e;
         2868: data_out <= 8'h60;
         2869: data_out <= 8'h81;
         2870: data_out <= 8'h9e;
         2871: data_out <= 8'h26;
         2872: data_out <= 8'h03;
         2873: data_out <= 8'h7e;
         2874: data_out <= 8'h0e;
         2875: data_out <= 8'hb9;
         2876: data_out <= 8'h80;
         2877: data_out <= 8'had;
         2878: data_out <= 8'h24;
         2879: data_out <= 8'h30;
         2880: data_out <= 8'h8d;
         2881: data_out <= 8'h06;
         2882: data_out <= 8'hbd;
         2883: data_out <= 8'h0a;
         2884: data_out <= 8'h27;
         2885: data_out <= 8'hc6;
         2886: data_out <= 8'h29;
         2887: data_out <= 8'h8c;
         2888: data_out <= 8'hc6;
         2889: data_out <= 8'h28;
         2890: data_out <= 8'h8c;
         2891: data_out <= 8'hc6;
         2892: data_out <= 8'h2c;
         2893: data_out <= 8'hde;
         2894: data_out <= 8'hc8;
         2895: data_out <= 8'ha6;
         2896: data_out <= 8'h00;
         2897: data_out <= 8'h11;
         2898: data_out <= 8'h26;
         2899: data_out <= 8'h03;
         2900: data_out <= 8'h7e;
         2901: data_out <= 8'h00;
         2902: data_out <= 8'hbf;
         2903: data_out <= 8'hc6;
         2904: data_out <= 8'h02;
         2905: data_out <= 8'h7e;
         2906: data_out <= 8'h03;
         2907: data_out <= 8'h21;
         2908: data_out <= 8'h86;
         2909: data_out <= 8'h7d;
         2910: data_out <= 8'hbd;
         2911: data_out <= 8'h0a;
         2912: data_out <= 8'h2e;
         2913: data_out <= 8'h7e;
         2914: data_out <= 8'h18;
         2915: data_out <= 8'h91;
         2916: data_out <= 8'hbd;
         2917: data_out <= 8'h0c;
         2918: data_out <= 8'h37;
         2919: data_out <= 8'hdf;
         2920: data_out <= 8'hb1;
         2921: data_out <= 8'h96;
         2922: data_out <= 8'h5c;
         2923: data_out <= 8'h26;
         2924: data_out <= 8'h8b;
         2925: data_out <= 8'h7e;
         2926: data_out <= 8'h15;
         2927: data_out <= 8'h8e;
         2928: data_out <= 8'h16;
         2929: data_out <= 8'h58;
         2930: data_out <= 8'h8d;
         2931: data_out <= 8'he0;
         2932: data_out <= 8'h37;
         2933: data_out <= 8'hc1;
         2934: data_out <= 8'h27;
         2935: data_out <= 8'h25;
         2936: data_out <= 8'h1a;
         2937: data_out <= 8'h8d;
         2938: data_out <= 8'hcd;
         2939: data_out <= 8'hbd;
         2940: data_out <= 8'h0a;
         2941: data_out <= 8'h27;
         2942: data_out <= 8'h8d;
         2943: data_out <= 8'hcb;
         2944: data_out <= 8'hbd;
         2945: data_out <= 8'h0a;
         2946: data_out <= 8'h1c;
         2947: data_out <= 8'h32;
         2948: data_out <= 8'hd6;
         2949: data_out <= 8'hb2;
         2950: data_out <= 8'h37;
         2951: data_out <= 8'hd6;
         2952: data_out <= 8'hb1;
         2953: data_out <= 8'h37;
         2954: data_out <= 8'h36;
         2955: data_out <= 8'hbd;
         2956: data_out <= 8'h11;
         2957: data_out <= 8'h6a;
         2958: data_out <= 8'h32;
         2959: data_out <= 8'h37;
         2960: data_out <= 8'h16;
         2961: data_out <= 8'h20;
         2962: data_out <= 8'h03;
         2963: data_out <= 8'h8d;
         2964: data_out <= 8'hab;
         2965: data_out <= 8'h33;
         2966: data_out <= 8'hce;
         2967: data_out <= 8'h01;
         2968: data_out <= 8'h19;
         2969: data_out <= 8'hbd;
         2970: data_out <= 8'h03;
         2971: data_out <= 8'h11;
         2972: data_out <= 8'hee;
         2973: data_out <= 8'h00;
         2974: data_out <= 8'had;
         2975: data_out <= 8'h00;
         2976: data_out <= 8'h7e;
         2977: data_out <= 8'h0a;
         2978: data_out <= 8'h1b;
         2979: data_out <= 8'h86;
         2980: data_out <= 8'h4f;
         2981: data_out <= 8'h97;
         2982: data_out <= 8'h5a;
         2983: data_out <= 8'hbd;
         2984: data_out <= 8'h0c;
         2985: data_out <= 8'hf1;
         2986: data_out <= 8'hde;
         2987: data_out <= 8'hb1;
         2988: data_out <= 8'hdf;
         2989: data_out <= 8'h58;
         2990: data_out <= 8'hbd;
         2991: data_out <= 8'h15;
         2992: data_out <= 8'hbf;
         2993: data_out <= 8'hbd;
         2994: data_out <= 8'h0c;
         2995: data_out <= 8'hf1;
         2996: data_out <= 8'h96;
         2997: data_out <= 8'h58;
         2998: data_out <= 8'hd6;
         2999: data_out <= 8'h59;
         3000: data_out <= 8'h7d;
         3001: data_out <= 8'h00;
         3002: data_out <= 8'h5a;
         3003: data_out <= 8'h26;
         3004: data_out <= 8'h06;
         3005: data_out <= 8'h94;
         3006: data_out <= 8'hb1;
         3007: data_out <= 8'hd4;
         3008: data_out <= 8'hb2;
         3009: data_out <= 8'h20;
         3010: data_out <= 8'h04;
         3011: data_out <= 8'h9a;
         3012: data_out <= 8'hb1;
         3013: data_out <= 8'hda;
         3014: data_out <= 8'hb2;
         3015: data_out <= 8'h7e;
         3016: data_out <= 8'h0e;
         3017: data_out <= 8'h60;
         3018: data_out <= 8'hbd;
         3019: data_out <= 8'h0a;
         3020: data_out <= 8'h1d;
         3021: data_out <= 8'h26;
         3022: data_out <= 8'h10;
         3023: data_out <= 8'h96;
         3024: data_out <= 8'hba;
         3025: data_out <= 8'h8a;
         3026: data_out <= 8'h7f;
         3027: data_out <= 8'h94;
         3028: data_out <= 8'hb7;
         3029: data_out <= 8'h97;
         3030: data_out <= 8'hb7;
         3031: data_out <= 8'hce;
         3032: data_out <= 8'h00;
         3033: data_out <= 8'hb6;
         3034: data_out <= 8'hbd;
         3035: data_out <= 8'h16;
         3036: data_out <= 8'h04;
         3037: data_out <= 8'h20;
         3038: data_out <= 8'h40;
         3039: data_out <= 8'h7f;
         3040: data_out <= 8'h00;
         3041: data_out <= 8'h5c;
         3042: data_out <= 8'h7a;
         3043: data_out <= 8'h00;
         3044: data_out <= 8'ha2;
         3045: data_out <= 8'hbd;
         3046: data_out <= 8'h10;
         3047: data_out <= 8'ha9;
         3048: data_out <= 8'hd7;
         3049: data_out <= 8'haf;
         3050: data_out <= 8'hdf;
         3051: data_out <= 8'hb1;
         3052: data_out <= 8'hde;
         3053: data_out <= 8'hb8;
         3054: data_out <= 8'hbd;
         3055: data_out <= 8'h10;
         3056: data_out <= 8'hab;
         3057: data_out <= 8'h96;
         3058: data_out <= 8'haf;
         3059: data_out <= 8'h10;
         3060: data_out <= 8'h27;
         3061: data_out <= 8'h07;
         3062: data_out <= 8'h86;
         3063: data_out <= 8'h01;
         3064: data_out <= 8'h24;
         3065: data_out <= 8'h03;
         3066: data_out <= 8'hd6;
         3067: data_out <= 8'haf;
         3068: data_out <= 8'h40;
         3069: data_out <= 8'h97;
         3070: data_out <= 8'hb3;
         3071: data_out <= 8'h07;
         3072: data_out <= 8'h36;
         3073: data_out <= 8'h9f;
         3074: data_out <= 8'h78;
         3075: data_out <= 8'h0f;
         3076: data_out <= 8'h35;
         3077: data_out <= 8'hde;
         3078: data_out <= 8'hb1;
         3079: data_out <= 8'h5c;
         3080: data_out <= 8'h09;
         3081: data_out <= 8'h5a;
         3082: data_out <= 8'h26;
         3083: data_out <= 8'h04;
         3084: data_out <= 8'hd6;
         3085: data_out <= 8'hb3;
         3086: data_out <= 8'h20;
         3087: data_out <= 8'h0b;
         3088: data_out <= 8'h32;
         3089: data_out <= 8'h08;
         3090: data_out <= 8'ha1;
         3091: data_out <= 8'h00;
         3092: data_out <= 8'h27;
         3093: data_out <= 8'hf3;
         3094: data_out <= 8'hc6;
         3095: data_out <= 8'hff;
         3096: data_out <= 8'h24;
         3097: data_out <= 8'h01;
         3098: data_out <= 8'h50;
         3099: data_out <= 8'h9e;
         3100: data_out <= 8'h78;
         3101: data_out <= 8'h32;
         3102: data_out <= 8'h06;
         3103: data_out <= 8'hcb;
         3104: data_out <= 8'h01;
         3105: data_out <= 8'h59;
         3106: data_out <= 8'hd4;
         3107: data_out <= 8'h60;
         3108: data_out <= 8'h27;
         3109: data_out <= 8'h02;
         3110: data_out <= 8'hc6;
         3111: data_out <= 8'hff;
         3112: data_out <= 8'h7e;
         3113: data_out <= 8'h15;
         3114: data_out <= 8'he8;
         3115: data_out <= 8'hbd;
         3116: data_out <= 8'h0b;
         3117: data_out <= 8'h4b;
         3118: data_out <= 8'h16;
         3119: data_out <= 8'h8d;
         3120: data_out <= 8'h0a;
         3121: data_out <= 8'hbd;
         3122: data_out <= 8'h00;
         3123: data_out <= 8'hc7;
         3124: data_out <= 8'h26;
         3125: data_out <= 8'hf5;
         3126: data_out <= 8'h39;
         3127: data_out <= 8'h5f;
         3128: data_out <= 8'hbd;
         3129: data_out <= 8'h00;
         3130: data_out <= 8'hc7;
         3131: data_out <= 8'hd7;
         3132: data_out <= 8'h5b;
         3133: data_out <= 8'h97;
         3134: data_out <= 8'h9a;
         3135: data_out <= 8'hbd;
         3136: data_out <= 8'h00;
         3137: data_out <= 8'hc7;
         3138: data_out <= 8'h8d;
         3139: data_out <= 8'h57;
         3140: data_out <= 8'h24;
         3141: data_out <= 8'h03;
         3142: data_out <= 8'h7e;
         3143: data_out <= 8'h0b;
         3144: data_out <= 8'h57;
         3145: data_out <= 8'h5f;
         3146: data_out <= 8'hd7;
         3147: data_out <= 8'h5c;
         3148: data_out <= 8'hbd;
         3149: data_out <= 8'h00;
         3150: data_out <= 8'hbf;
         3151: data_out <= 8'h25;
         3152: data_out <= 8'h04;
         3153: data_out <= 8'h8d;
         3154: data_out <= 8'h48;
         3155: data_out <= 8'h25;
         3156: data_out <= 8'h0a;
         3157: data_out <= 8'h16;
         3158: data_out <= 8'hbd;
         3159: data_out <= 8'h00;
         3160: data_out <= 8'hbf;
         3161: data_out <= 8'h25;
         3162: data_out <= 8'hfb;
         3163: data_out <= 8'h8d;
         3164: data_out <= 8'h3e;
         3165: data_out <= 8'h24;
         3166: data_out <= 8'hf7;
         3167: data_out <= 8'h81;
         3168: data_out <= 8'h24;
         3169: data_out <= 8'h26;
         3170: data_out <= 8'h08;
         3171: data_out <= 8'h73;
         3172: data_out <= 8'h00;
         3173: data_out <= 8'h5c;
         3174: data_out <= 8'hcb;
         3175: data_out <= 8'h80;
         3176: data_out <= 8'hbd;
         3177: data_out <= 8'h00;
         3178: data_out <= 8'hbf;
         3179: data_out <= 8'hd7;
         3180: data_out <= 8'h9b;
         3181: data_out <= 8'hd6;
         3182: data_out <= 8'h5e;
         3183: data_out <= 8'h5a;
         3184: data_out <= 8'h26;
         3185: data_out <= 8'h03;
         3186: data_out <= 8'h7e;
         3187: data_out <= 8'h0d;
         3188: data_out <= 8'h3e;
         3189: data_out <= 8'h9b;
         3190: data_out <= 8'h5e;
         3191: data_out <= 8'h80;
         3192: data_out <= 8'h28;
         3193: data_out <= 8'h26;
         3194: data_out <= 8'h03;
         3195: data_out <= 8'h7e;
         3196: data_out <= 8'h0d;
         3197: data_out <= 8'h02;
         3198: data_out <= 8'h7f;
         3199: data_out <= 8'h00;
         3200: data_out <= 8'h5e;
         3201: data_out <= 8'hde;
         3202: data_out <= 8'h7c;
         3203: data_out <= 8'h96;
         3204: data_out <= 8'h9a;
         3205: data_out <= 8'hd6;
         3206: data_out <= 8'h9b;
         3207: data_out <= 8'h9c;
         3208: data_out <= 8'h7e;
         3209: data_out <= 8'h27;
         3210: data_out <= 8'h19;
         3211: data_out <= 8'ha1;
         3212: data_out <= 8'h00;
         3213: data_out <= 8'h26;
         3214: data_out <= 8'h04;
         3215: data_out <= 8'he1;
         3216: data_out <= 8'h01;
         3217: data_out <= 8'h27;
         3218: data_out <= 8'h48;
         3219: data_out <= 8'h08;
         3220: data_out <= 8'h08;
         3221: data_out <= 8'h08;
         3222: data_out <= 8'h08;
         3223: data_out <= 8'h08;
         3224: data_out <= 8'h08;
         3225: data_out <= 8'h20;
         3226: data_out <= 8'hec;
         3227: data_out <= 8'h81;
         3228: data_out <= 8'h41;
         3229: data_out <= 8'h25;
         3230: data_out <= 8'h04;
         3231: data_out <= 8'h80;
         3232: data_out <= 8'h5b;
         3233: data_out <= 8'h80;
         3234: data_out <= 8'ha5;
         3235: data_out <= 8'h39;
         3236: data_out <= 8'h32;
         3237: data_out <= 8'h36;
         3238: data_out <= 8'h81;
         3239: data_out <= 8'h0b;
         3240: data_out <= 8'h26;
         3241: data_out <= 8'h04;
         3242: data_out <= 8'hce;
         3243: data_out <= 8'h0d;
         3244: data_out <= 8'h1e;
         3245: data_out <= 8'h39;
         3246: data_out <= 8'hde;
         3247: data_out <= 8'h80;
         3248: data_out <= 8'hdf;
         3249: data_out <= 8'ha5;
         3250: data_out <= 8'hc6;
         3251: data_out <= 8'h06;
         3252: data_out <= 8'hbd;
         3253: data_out <= 8'h03;
         3254: data_out <= 8'h11;
         3255: data_out <= 8'hdf;
         3256: data_out <= 8'ha3;
         3257: data_out <= 8'hde;
         3258: data_out <= 8'h7e;
         3259: data_out <= 8'hdf;
         3260: data_out <= 8'ha9;
         3261: data_out <= 8'hbd;
         3262: data_out <= 8'h02;
         3263: data_out <= 8'hdc;
         3264: data_out <= 8'hde;
         3265: data_out <= 8'ha3;
         3266: data_out <= 8'hdf;
         3267: data_out <= 8'h80;
         3268: data_out <= 8'hde;
         3269: data_out <= 8'ha7;
         3270: data_out <= 8'hdf;
         3271: data_out <= 8'h7e;
         3272: data_out <= 8'hde;
         3273: data_out <= 8'ha9;
         3274: data_out <= 8'h96;
         3275: data_out <= 8'h9a;
         3276: data_out <= 8'hd6;
         3277: data_out <= 8'h9b;
         3278: data_out <= 8'ha7;
         3279: data_out <= 8'h00;
         3280: data_out <= 8'he7;
         3281: data_out <= 8'h01;
         3282: data_out <= 8'h4f;
         3283: data_out <= 8'ha7;
         3284: data_out <= 8'h02;
         3285: data_out <= 8'ha7;
         3286: data_out <= 8'h03;
         3287: data_out <= 8'ha7;
         3288: data_out <= 8'h04;
         3289: data_out <= 8'ha7;
         3290: data_out <= 8'h05;
         3291: data_out <= 8'h08;
         3292: data_out <= 8'h08;
         3293: data_out <= 8'hdf;
         3294: data_out <= 8'h9c;
         3295: data_out <= 8'h39;
         3296: data_out <= 8'h90;
         3297: data_out <= 8'h80;
         3298: data_out <= 8'h00;
         3299: data_out <= 8'h00;
         3300: data_out <= 8'hbd;
         3301: data_out <= 8'h00;
         3302: data_out <= 8'hbf;
         3303: data_out <= 8'hbd;
         3304: data_out <= 8'h0a;
         3305: data_out <= 8'h19;
         3306: data_out <= 8'h96;
         3307: data_out <= 8'hb3;
         3308: data_out <= 8'h2a;
         3309: data_out <= 8'h03;
         3310: data_out <= 8'h7e;
         3311: data_out <= 8'h0d;
         3312: data_out <= 8'h71;
         3313: data_out <= 8'h96;
         3314: data_out <= 8'haf;
         3315: data_out <= 8'h81;
         3316: data_out <= 8'h90;
         3317: data_out <= 8'h25;
         3318: data_out <= 8'h08;
         3319: data_out <= 8'hce;
         3320: data_out <= 8'h0c;
         3321: data_out <= 8'he0;
         3322: data_out <= 8'hbd;
         3323: data_out <= 8'h16;
         3324: data_out <= 8'h04;
         3325: data_out <= 8'h26;
         3326: data_out <= 8'h72;
         3327: data_out <= 8'h7e;
         3328: data_out <= 8'h16;
         3329: data_out <= 8'h30;
         3330: data_out <= 8'h96;
         3331: data_out <= 8'h5b;
         3332: data_out <= 8'h36;
         3333: data_out <= 8'h96;
         3334: data_out <= 8'h5c;
         3335: data_out <= 8'h36;
         3336: data_out <= 8'h5f;
         3337: data_out <= 8'h37;
         3338: data_out <= 8'hd6;
         3339: data_out <= 8'h9b;
         3340: data_out <= 8'h37;
         3341: data_out <= 8'hd6;
         3342: data_out <= 8'h9a;
         3343: data_out <= 8'h37;
         3344: data_out <= 8'h8d;
         3345: data_out <= 8'hd2;
         3346: data_out <= 8'h33;
         3347: data_out <= 8'hd7;
         3348: data_out <= 8'h9a;
         3349: data_out <= 8'h33;
         3350: data_out <= 8'hd7;
         3351: data_out <= 8'h9b;
         3352: data_out <= 8'h33;
         3353: data_out <= 8'h30;
         3354: data_out <= 8'ha6;
         3355: data_out <= 8'h01;
         3356: data_out <= 8'h36;
         3357: data_out <= 8'ha6;
         3358: data_out <= 8'h00;
         3359: data_out <= 8'h36;
         3360: data_out <= 8'h96;
         3361: data_out <= 8'hb1;
         3362: data_out <= 8'ha7;
         3363: data_out <= 8'h00;
         3364: data_out <= 8'h96;
         3365: data_out <= 8'hb2;
         3366: data_out <= 8'ha7;
         3367: data_out <= 8'h01;
         3368: data_out <= 8'h5c;
         3369: data_out <= 8'hbd;
         3370: data_out <= 8'h00;
         3371: data_out <= 8'hc7;
         3372: data_out <= 8'h81;
         3373: data_out <= 8'h2c;
         3374: data_out <= 8'h27;
         3375: data_out <= 8'hd9;
         3376: data_out <= 8'hd7;
         3377: data_out <= 8'h5a;
         3378: data_out <= 8'hbd;
         3379: data_out <= 8'h0b;
         3380: data_out <= 8'h45;
         3381: data_out <= 8'h32;
         3382: data_out <= 8'h97;
         3383: data_out <= 8'h5c;
         3384: data_out <= 8'h32;
         3385: data_out <= 8'h97;
         3386: data_out <= 8'h5b;
         3387: data_out <= 8'hc6;
         3388: data_out <= 8'hff;
         3389: data_out <= 8'h86;
         3390: data_out <= 8'h5f;
         3391: data_out <= 8'h37;
         3392: data_out <= 8'hde;
         3393: data_out <= 8'h7e;
         3394: data_out <= 8'h9c;
         3395: data_out <= 8'h80;
         3396: data_out <= 8'h27;
         3397: data_out <= 8'h30;
         3398: data_out <= 8'h96;
         3399: data_out <= 8'h9a;
         3400: data_out <= 8'ha1;
         3401: data_out <= 8'h00;
         3402: data_out <= 8'h26;
         3403: data_out <= 8'h06;
         3404: data_out <= 8'h96;
         3405: data_out <= 8'h9b;
         3406: data_out <= 8'ha1;
         3407: data_out <= 8'h01;
         3408: data_out <= 8'h27;
         3409: data_out <= 8'h09;
         3410: data_out <= 8'ha6;
         3411: data_out <= 8'h02;
         3412: data_out <= 8'he6;
         3413: data_out <= 8'h03;
         3414: data_out <= 8'hbd;
         3415: data_out <= 8'h03;
         3416: data_out <= 8'h12;
         3417: data_out <= 8'h20;
         3418: data_out <= 8'he7;
         3419: data_out <= 8'hc6;
         3420: data_out <= 8'h12;
         3421: data_out <= 8'h32;
         3422: data_out <= 8'h4d;
         3423: data_out <= 8'h26;
         3424: data_out <= 8'h03;
         3425: data_out <= 8'h7e;
         3426: data_out <= 8'h12;
         3427: data_out <= 8'hb4;
         3428: data_out <= 8'h96;
         3429: data_out <= 8'h5b;
         3430: data_out <= 8'h26;
         3431: data_out <= 8'h0b;
         3432: data_out <= 8'hd6;
         3433: data_out <= 8'h5a;
         3434: data_out <= 8'he1;
         3435: data_out <= 8'h04;
         3436: data_out <= 8'h27;
         3437: data_out <= 8'h6e;
         3438: data_out <= 8'hc6;
         3439: data_out <= 8'h10;
         3440: data_out <= 8'h8c;
         3441: data_out <= 8'hc6;
         3442: data_out <= 8'h08;
         3443: data_out <= 8'h7e;
         3444: data_out <= 8'h03;
         3445: data_out <= 8'h21;
         3446: data_out <= 8'h32;
         3447: data_out <= 8'h4d;
         3448: data_out <= 8'h26;
         3449: data_out <= 8'h03;
         3450: data_out <= 8'h7e;
         3451: data_out <= 8'h0b;
         3452: data_out <= 8'h57;
         3453: data_out <= 8'h86;
         3454: data_out <= 8'h04;
         3455: data_out <= 8'h97;
         3456: data_out <= 8'hbe;
         3457: data_out <= 8'h7f;
         3458: data_out <= 8'h00;
         3459: data_out <= 8'hbd;
         3460: data_out <= 8'h96;
         3461: data_out <= 8'h9a;
         3462: data_out <= 8'ha7;
         3463: data_out <= 8'h00;
         3464: data_out <= 8'h96;
         3465: data_out <= 8'h9b;
         3466: data_out <= 8'ha7;
         3467: data_out <= 8'h01;
         3468: data_out <= 8'hd6;
         3469: data_out <= 8'h5a;
         3470: data_out <= 8'he7;
         3471: data_out <= 8'h04;
         3472: data_out <= 8'hbd;
         3473: data_out <= 8'h02;
         3474: data_out <= 8'hf8;
         3475: data_out <= 8'hdf;
         3476: data_out <= 8'ha3;
         3477: data_out <= 8'hc6;
         3478: data_out <= 8'h0b;
         3479: data_out <= 8'h4f;
         3480: data_out <= 8'h7d;
         3481: data_out <= 8'h00;
         3482: data_out <= 8'h5b;
         3483: data_out <= 8'h27;
         3484: data_out <= 8'h06;
         3485: data_out <= 8'h32;
         3486: data_out <= 8'h33;
         3487: data_out <= 8'hcb;
         3488: data_out <= 8'h01;
         3489: data_out <= 8'h89;
         3490: data_out <= 8'h00;
         3491: data_out <= 8'ha7;
         3492: data_out <= 8'h05;
         3493: data_out <= 8'he7;
         3494: data_out <= 8'h06;
         3495: data_out <= 8'h8d;
         3496: data_out <= 8'h6f;
         3497: data_out <= 8'h97;
         3498: data_out <= 8'hbd;
         3499: data_out <= 8'hd7;
         3500: data_out <= 8'hbe;
         3501: data_out <= 8'h08;
         3502: data_out <= 8'h08;
         3503: data_out <= 8'h7a;
         3504: data_out <= 8'h00;
         3505: data_out <= 8'h5a;
         3506: data_out <= 8'h26;
         3507: data_out <= 8'he1;
         3508: data_out <= 8'hbd;
         3509: data_out <= 8'h03;
         3510: data_out <= 8'h12;
         3511: data_out <= 8'h25;
         3512: data_out <= 8'hb5;
         3513: data_out <= 8'hbd;
         3514: data_out <= 8'h02;
         3515: data_out <= 8'hfe;
         3516: data_out <= 8'hc0;
         3517: data_out <= 8'h21;
         3518: data_out <= 8'h82;
         3519: data_out <= 8'h00;
         3520: data_out <= 8'h97;
         3521: data_out <= 8'h80;
         3522: data_out <= 8'hd7;
         3523: data_out <= 8'h81;
         3524: data_out <= 8'h4f;
         3525: data_out <= 8'h09;
         3526: data_out <= 8'ha7;
         3527: data_out <= 8'h05;
         3528: data_out <= 8'h9c;
         3529: data_out <= 8'h71;
         3530: data_out <= 8'h26;
         3531: data_out <= 8'hf9;
         3532: data_out <= 8'hde;
         3533: data_out <= 8'ha3;
         3534: data_out <= 8'h96;
         3535: data_out <= 8'h80;
         3536: data_out <= 8'hd0;
         3537: data_out <= 8'ha4;
         3538: data_out <= 8'he7;
         3539: data_out <= 8'h03;
         3540: data_out <= 8'h92;
         3541: data_out <= 8'ha3;
         3542: data_out <= 8'ha7;
         3543: data_out <= 8'h02;
         3544: data_out <= 8'h96;
         3545: data_out <= 8'h5b;
         3546: data_out <= 8'h26;
         3547: data_out <= 8'h3b;
         3548: data_out <= 8'he6;
         3549: data_out <= 8'h04;
         3550: data_out <= 8'hd7;
         3551: data_out <= 8'h5a;
         3552: data_out <= 8'h4f;
         3553: data_out <= 8'h5f;
         3554: data_out <= 8'h97;
         3555: data_out <= 8'hbd;
         3556: data_out <= 8'hd7;
         3557: data_out <= 8'hbe;
         3558: data_out <= 8'h32;
         3559: data_out <= 8'h97;
         3560: data_out <= 8'hb1;
         3561: data_out <= 8'h33;
         3562: data_out <= 8'hd7;
         3563: data_out <= 8'hb2;
         3564: data_out <= 8'ha1;
         3565: data_out <= 8'h05;
         3566: data_out <= 8'h25;
         3567: data_out <= 8'h06;
         3568: data_out <= 8'h22;
         3569: data_out <= 8'h4c;
         3570: data_out <= 8'he1;
         3571: data_out <= 8'h06;
         3572: data_out <= 8'h24;
         3573: data_out <= 8'h48;
         3574: data_out <= 8'h96;
         3575: data_out <= 8'hbe;
         3576: data_out <= 8'h9a;
         3577: data_out <= 8'hbd;
         3578: data_out <= 8'h0c;
         3579: data_out <= 8'h27;
         3580: data_out <= 8'h04;
         3581: data_out <= 8'h8d;
         3582: data_out <= 8'h19;
         3583: data_out <= 8'hdb;
         3584: data_out <= 8'hb2;
         3585: data_out <= 8'h99;
         3586: data_out <= 8'hb1;
         3587: data_out <= 8'h08;
         3588: data_out <= 8'h08;
         3589: data_out <= 8'h7a;
         3590: data_out <= 8'h00;
         3591: data_out <= 8'h5a;
         3592: data_out <= 8'h26;
         3593: data_out <= 8'hd8;
         3594: data_out <= 8'h58;
         3595: data_out <= 8'h49;
         3596: data_out <= 8'h58;
         3597: data_out <= 8'h49;
         3598: data_out <= 8'hcb;
         3599: data_out <= 8'h05;
         3600: data_out <= 8'h89;
         3601: data_out <= 8'h00;
         3602: data_out <= 8'hbd;
         3603: data_out <= 8'h03;
         3604: data_out <= 8'h12;
         3605: data_out <= 8'hdf;
         3606: data_out <= 8'h9c;
         3607: data_out <= 8'h39;
         3608: data_out <= 8'h86;
         3609: data_out <= 8'h10;
         3610: data_out <= 8'h97;
         3611: data_out <= 8'ha7;
         3612: data_out <= 8'ha6;
         3613: data_out <= 8'h05;
         3614: data_out <= 8'h97;
         3615: data_out <= 8'h78;
         3616: data_out <= 8'ha6;
         3617: data_out <= 8'h06;
         3618: data_out <= 8'h97;
         3619: data_out <= 8'h79;
         3620: data_out <= 8'h4f;
         3621: data_out <= 8'h5f;
         3622: data_out <= 8'h58;
         3623: data_out <= 8'h49;
         3624: data_out <= 8'h25;
         3625: data_out <= 8'h14;
         3626: data_out <= 8'h78;
         3627: data_out <= 8'h00;
         3628: data_out <= 8'hbe;
         3629: data_out <= 8'h79;
         3630: data_out <= 8'h00;
         3631: data_out <= 8'hbd;
         3632: data_out <= 8'h24;
         3633: data_out <= 8'h06;
         3634: data_out <= 8'hdb;
         3635: data_out <= 8'h79;
         3636: data_out <= 8'h99;
         3637: data_out <= 8'h78;
         3638: data_out <= 8'h25;
         3639: data_out <= 8'h06;
         3640: data_out <= 8'h7a;
         3641: data_out <= 8'h00;
         3642: data_out <= 8'ha7;
         3643: data_out <= 8'h26;
         3644: data_out <= 8'he9;
         3645: data_out <= 8'h39;
         3646: data_out <= 8'h7e;
         3647: data_out <= 8'h0d;
         3648: data_out <= 8'h6e;
         3649: data_out <= 8'h9f;
         3650: data_out <= 8'h78;
         3651: data_out <= 8'h96;
         3652: data_out <= 8'h78;
         3653: data_out <= 8'hd6;
         3654: data_out <= 8'h79;
         3655: data_out <= 8'hce;
         3656: data_out <= 8'h00;
         3657: data_out <= 8'h80;
         3658: data_out <= 8'h7d;
         3659: data_out <= 8'h00;
         3660: data_out <= 8'h5c;
         3661: data_out <= 8'h27;
         3662: data_out <= 8'h0d;
         3663: data_out <= 8'hbd;
         3664: data_out <= 8'h10;
         3665: data_out <= 8'ha9;
         3666: data_out <= 8'hbd;
         3667: data_out <= 8'h0f;
         3668: data_out <= 8'hb2;
         3669: data_out <= 8'hce;
         3670: data_out <= 8'h00;
         3671: data_out <= 8'h82;
         3672: data_out <= 8'h96;
         3673: data_out <= 8'h84;
         3674: data_out <= 8'hd6;
         3675: data_out <= 8'h85;
         3676: data_out <= 8'he0;
         3677: data_out <= 8'h01;
         3678: data_out <= 8'ha2;
         3679: data_out <= 8'h00;
         3680: data_out <= 8'h7f;
         3681: data_out <= 8'h00;
         3682: data_out <= 8'h5c;
         3683: data_out <= 8'h97;
         3684: data_out <= 8'hb0;
         3685: data_out <= 8'hd7;
         3686: data_out <= 8'hb1;
         3687: data_out <= 8'hc6;
         3688: data_out <= 8'h90;
         3689: data_out <= 8'h7e;
         3690: data_out <= 8'h15;
         3691: data_out <= 8'hef;
         3692: data_out <= 8'hd6;
         3693: data_out <= 8'h0b;
         3694: data_out <= 8'h4f;
         3695: data_out <= 8'h20;
         3696: data_out <= 8'hef;
         3697: data_out <= 8'hde;
         3698: data_out <= 8'h8a;
         3699: data_out <= 8'h08;
         3700: data_out <= 8'h26;
         3701: data_out <= 8'ha1;
         3702: data_out <= 8'hc6;
         3703: data_out <= 8'h16;
         3704: data_out <= 8'h7e;
         3705: data_out <= 8'h03;
         3706: data_out <= 8'h21;
         3707: data_out <= 8'h8d;
         3708: data_out <= 8'h29;
         3709: data_out <= 8'h8d;
         3710: data_out <= 8'hf2;
         3711: data_out <= 8'hbd;
         3712: data_out <= 8'h0b;
         3713: data_out <= 8'h48;
         3714: data_out <= 8'hc6;
         3715: data_out <= 8'h80;
         3716: data_out <= 8'hd7;
         3717: data_out <= 8'h5e;
         3718: data_out <= 8'hbd;
         3719: data_out <= 8'h0c;
         3720: data_out <= 8'h37;
         3721: data_out <= 8'h8d;
         3722: data_out <= 8'h2b;
         3723: data_out <= 8'hbd;
         3724: data_out <= 8'h0b;
         3725: data_out <= 8'h45;
         3726: data_out <= 8'hc6;
         3727: data_out <= 8'hab;
         3728: data_out <= 8'hbd;
         3729: data_out <= 8'h0b;
         3730: data_out <= 8'h4d;
         3731: data_out <= 8'hde;
         3732: data_out <= 8'hab;
         3733: data_out <= 8'h96;
         3734: data_out <= 8'hc8;
         3735: data_out <= 8'hd6;
         3736: data_out <= 8'hc9;
         3737: data_out <= 8'ha7;
         3738: data_out <= 8'h00;
         3739: data_out <= 8'he7;
         3740: data_out <= 8'h01;
         3741: data_out <= 8'h96;
         3742: data_out <= 8'h9c;
         3743: data_out <= 8'hd6;
         3744: data_out <= 8'h9d;
         3745: data_out <= 8'h8d;
         3746: data_out <= 8'h75;
         3747: data_out <= 8'h7e;
         3748: data_out <= 8'h07;
         3749: data_out <= 8'h14;
         3750: data_out <= 8'hc6;
         3751: data_out <= 8'h9e;
         3752: data_out <= 8'hbd;
         3753: data_out <= 8'h0b;
         3754: data_out <= 8'h4d;
         3755: data_out <= 8'hc6;
         3756: data_out <= 8'h80;
         3757: data_out <= 8'hd7;
         3758: data_out <= 8'h5e;
         3759: data_out <= 8'h8a;
         3760: data_out <= 8'h80;
         3761: data_out <= 8'hbd;
         3762: data_out <= 8'h0c;
         3763: data_out <= 8'h3d;
         3764: data_out <= 8'hdf;
         3765: data_out <= 8'hab;
         3766: data_out <= 8'h7e;
         3767: data_out <= 8'h0a;
         3768: data_out <= 8'h1b;
         3769: data_out <= 8'h8d;
         3770: data_out <= 8'heb;
         3771: data_out <= 8'hd6;
         3772: data_out <= 8'hac;
         3773: data_out <= 8'h37;
         3774: data_out <= 8'hd6;
         3775: data_out <= 8'hab;
         3776: data_out <= 8'h37;
         3777: data_out <= 8'hbd;
         3778: data_out <= 8'h0b;
         3779: data_out <= 8'h40;
         3780: data_out <= 8'h8d;
         3781: data_out <= 8'hf0;
         3782: data_out <= 8'h33;
         3783: data_out <= 8'hd7;
         3784: data_out <= 8'hab;
         3785: data_out <= 8'h33;
         3786: data_out <= 8'hd7;
         3787: data_out <= 8'hac;
         3788: data_out <= 8'hde;
         3789: data_out <= 8'hab;
         3790: data_out <= 8'hc6;
         3791: data_out <= 8'h22;
         3792: data_out <= 8'hee;
         3793: data_out <= 8'h02;
         3794: data_out <= 8'h27;
         3795: data_out <= 8'ha4;
         3796: data_out <= 8'hdf;
         3797: data_out <= 8'h9c;
         3798: data_out <= 8'ha6;
         3799: data_out <= 8'h03;
         3800: data_out <= 8'h36;
         3801: data_out <= 8'ha6;
         3802: data_out <= 8'h02;
         3803: data_out <= 8'h36;
         3804: data_out <= 8'ha6;
         3805: data_out <= 8'h01;
         3806: data_out <= 8'h36;
         3807: data_out <= 8'ha6;
         3808: data_out <= 8'h00;
         3809: data_out <= 8'h36;
         3810: data_out <= 8'hbd;
         3811: data_out <= 8'h15;
         3812: data_out <= 8'haa;
         3813: data_out <= 8'hde;
         3814: data_out <= 8'hab;
         3815: data_out <= 8'hd6;
         3816: data_out <= 8'hc9;
         3817: data_out <= 8'h37;
         3818: data_out <= 8'hd6;
         3819: data_out <= 8'hc8;
         3820: data_out <= 8'h37;
         3821: data_out <= 8'hee;
         3822: data_out <= 8'h00;
         3823: data_out <= 8'hdf;
         3824: data_out <= 8'hc8;
         3825: data_out <= 8'hd6;
         3826: data_out <= 8'h9d;
         3827: data_out <= 8'h37;
         3828: data_out <= 8'hd6;
         3829: data_out <= 8'h9c;
         3830: data_out <= 8'h37;
         3831: data_out <= 8'hbd;
         3832: data_out <= 8'h0a;
         3833: data_out <= 8'h19;
         3834: data_out <= 8'h33;
         3835: data_out <= 8'hd7;
         3836: data_out <= 8'h9c;
         3837: data_out <= 8'h33;
         3838: data_out <= 8'hd7;
         3839: data_out <= 8'h9d;
         3840: data_out <= 8'hbd;
         3841: data_out <= 8'h00;
         3842: data_out <= 8'hc7;
         3843: data_out <= 8'h27;
         3844: data_out <= 8'h03;
         3845: data_out <= 8'h7e;
         3846: data_out <= 8'h0b;
         3847: data_out <= 8'h57;
         3848: data_out <= 8'h33;
         3849: data_out <= 8'hd7;
         3850: data_out <= 8'hc8;
         3851: data_out <= 8'h33;
         3852: data_out <= 8'hd7;
         3853: data_out <= 8'hc9;
         3854: data_out <= 8'hde;
         3855: data_out <= 8'h9c;
         3856: data_out <= 8'h32;
         3857: data_out <= 8'ha7;
         3858: data_out <= 8'h00;
         3859: data_out <= 8'h32;
         3860: data_out <= 8'ha7;
         3861: data_out <= 8'h01;
         3862: data_out <= 8'h32;
         3863: data_out <= 8'h33;
         3864: data_out <= 8'ha7;
         3865: data_out <= 8'h02;
         3866: data_out <= 8'he7;
         3867: data_out <= 8'h03;
         3868: data_out <= 8'h39;
         3869: data_out <= 8'hbd;
         3870: data_out <= 8'h0a;
         3871: data_out <= 8'h1b;
         3872: data_out <= 8'hce;
         3873: data_out <= 8'h00;
         3874: data_out <= 8'hff;
         3875: data_out <= 8'hbd;
         3876: data_out <= 8'h17;
         3877: data_out <= 8'h48;
         3878: data_out <= 8'h31;
         3879: data_out <= 8'h31;
         3880: data_out <= 8'hce;
         3881: data_out <= 8'h00;
         3882: data_out <= 8'hfe;
         3883: data_out <= 8'h20;
         3884: data_out <= 8'h0a;
         3885: data_out <= 8'hdf;
         3886: data_out <= 8'had;
         3887: data_out <= 8'h8d;
         3888: data_out <= 8'h53;
         3889: data_out <= 8'hdf;
         3890: data_out <= 8'hb1;
         3891: data_out <= 8'hd7;
         3892: data_out <= 8'haf;
         3893: data_out <= 8'h39;
         3894: data_out <= 8'h09;
         3895: data_out <= 8'h86;
         3896: data_out <= 8'h22;
         3897: data_out <= 8'h97;
         3898: data_out <= 8'h58;
         3899: data_out <= 8'h97;
         3900: data_out <= 8'h59;
         3901: data_out <= 8'h08;
         3902: data_out <= 8'hdf;
         3903: data_out <= 8'hbb;
         3904: data_out <= 8'hdf;
         3905: data_out <= 8'hb1;
         3906: data_out <= 8'hc6;
         3907: data_out <= 8'hff;
         3908: data_out <= 8'h5c;
         3909: data_out <= 8'ha6;
         3910: data_out <= 8'h00;
         3911: data_out <= 8'h27;
         3912: data_out <= 8'h0e;
         3913: data_out <= 8'h08;
         3914: data_out <= 8'h91;
         3915: data_out <= 8'h58;
         3916: data_out <= 8'h27;
         3917: data_out <= 8'h04;
         3918: data_out <= 8'h91;
         3919: data_out <= 8'h59;
         3920: data_out <= 8'h26;
         3921: data_out <= 8'hf2;
         3922: data_out <= 8'h81;
         3923: data_out <= 8'h22;
         3924: data_out <= 8'h27;
         3925: data_out <= 8'h01;
         3926: data_out <= 8'h09;
         3927: data_out <= 8'hdf;
         3928: data_out <= 8'hbd;
         3929: data_out <= 8'hd7;
         3930: data_out <= 8'haf;
         3931: data_out <= 8'h96;
         3932: data_out <= 8'hbb;
         3933: data_out <= 8'h26;
         3934: data_out <= 8'h07;
         3935: data_out <= 8'h8d;
         3936: data_out <= 8'hcc;
         3937: data_out <= 8'hde;
         3938: data_out <= 8'hbb;
         3939: data_out <= 8'hbd;
         3940: data_out <= 8'h10;
         3941: data_out <= 8'h8d;
         3942: data_out <= 8'hde;
         3943: data_out <= 8'h61;
         3944: data_out <= 8'h8c;
         3945: data_out <= 8'h00;
         3946: data_out <= 8'h71;
         3947: data_out <= 8'h26;
         3948: data_out <= 8'h05;
         3949: data_out <= 8'hc6;
         3950: data_out <= 8'h1e;
         3951: data_out <= 8'h7e;
         3952: data_out <= 8'h03;
         3953: data_out <= 8'h21;
         3954: data_out <= 8'hbd;
         3955: data_out <= 8'h15;
         3956: data_out <= 8'haa;
         3957: data_out <= 8'h86;
         3958: data_out <= 8'hff;
         3959: data_out <= 8'h97;
         3960: data_out <= 8'h5c;
         3961: data_out <= 8'hdf;
         3962: data_out <= 8'h63;
         3963: data_out <= 8'hdf;
         3964: data_out <= 8'hb1;
         3965: data_out <= 8'h08;
         3966: data_out <= 8'h08;
         3967: data_out <= 8'h08;
         3968: data_out <= 8'h08;
         3969: data_out <= 8'hdf;
         3970: data_out <= 8'h61;
         3971: data_out <= 8'h39;
         3972: data_out <= 8'h7f;
         3973: data_out <= 8'h00;
         3974: data_out <= 8'h5d;
         3975: data_out <= 8'h37;
         3976: data_out <= 8'h53;
         3977: data_out <= 8'h86;
         3978: data_out <= 8'hff;
         3979: data_out <= 8'hd9;
         3980: data_out <= 8'h85;
         3981: data_out <= 8'h99;
         3982: data_out <= 8'h84;
         3983: data_out <= 8'h91;
         3984: data_out <= 8'h82;
         3985: data_out <= 8'h25;
         3986: data_out <= 8'h11;
         3987: data_out <= 8'h22;
         3988: data_out <= 8'h04;
         3989: data_out <= 8'hd1;
         3990: data_out <= 8'h83;
         3991: data_out <= 8'h25;
         3992: data_out <= 8'h0b;
         3993: data_out <= 8'h97;
         3994: data_out <= 8'h84;
         3995: data_out <= 8'hd7;
         3996: data_out <= 8'h85;
         3997: data_out <= 8'hde;
         3998: data_out <= 8'h84;
         3999: data_out <= 8'h08;
         4000: data_out <= 8'hdf;
         4001: data_out <= 8'h86;
         4002: data_out <= 8'h33;
         4003: data_out <= 8'h39;
         4004: data_out <= 8'hc6;
         4005: data_out <= 8'h1a;
         4006: data_out <= 8'h96;
         4007: data_out <= 8'h5d;
         4008: data_out <= 8'h26;
         4009: data_out <= 8'hc5;
         4010: data_out <= 8'h8d;
         4011: data_out <= 8'h06;
         4012: data_out <= 8'h73;
         4013: data_out <= 8'h00;
         4014: data_out <= 8'h5d;
         4015: data_out <= 8'h33;
         4016: data_out <= 8'h20;
         4017: data_out <= 8'hd5;
         4018: data_out <= 8'hde;
         4019: data_out <= 8'h88;
         4020: data_out <= 8'hdf;
         4021: data_out <= 8'h84;
         4022: data_out <= 8'hce;
         4023: data_out <= 8'h00;
         4024: data_out <= 8'h00;
         4025: data_out <= 8'hdf;
         4026: data_out <= 8'hab;
         4027: data_out <= 8'hde;
         4028: data_out <= 8'h82;
         4029: data_out <= 8'hdf;
         4030: data_out <= 8'ha9;
         4031: data_out <= 8'hce;
         4032: data_out <= 8'h00;
         4033: data_out <= 8'h65;
         4034: data_out <= 8'h9c;
         4035: data_out <= 8'h61;
         4036: data_out <= 8'h27;
         4037: data_out <= 8'h04;
         4038: data_out <= 8'h8d;
         4039: data_out <= 8'h3b;
         4040: data_out <= 8'h20;
         4041: data_out <= 8'hf8;
         4042: data_out <= 8'hde;
         4043: data_out <= 8'h7c;
         4044: data_out <= 8'h9c;
         4045: data_out <= 8'h7e;
         4046: data_out <= 8'h27;
         4047: data_out <= 8'h04;
         4048: data_out <= 8'h8d;
         4049: data_out <= 8'h2b;
         4050: data_out <= 8'h20;
         4051: data_out <= 8'hf8;
         4052: data_out <= 8'hdf;
         4053: data_out <= 8'ha3;
         4054: data_out <= 8'hde;
         4055: data_out <= 8'ha3;
         4056: data_out <= 8'h9c;
         4057: data_out <= 8'h80;
         4058: data_out <= 8'h27;
         4059: data_out <= 8'h4e;
         4060: data_out <= 8'ha6;
         4061: data_out <= 8'h02;
         4062: data_out <= 8'he6;
         4063: data_out <= 8'h03;
         4064: data_out <= 8'hdb;
         4065: data_out <= 8'ha4;
         4066: data_out <= 8'h99;
         4067: data_out <= 8'ha3;
         4068: data_out <= 8'h97;
         4069: data_out <= 8'ha3;
         4070: data_out <= 8'hd7;
         4071: data_out <= 8'ha4;
         4072: data_out <= 8'ha6;
         4073: data_out <= 8'h01;
         4074: data_out <= 8'h2a;
         4075: data_out <= 8'hea;
         4076: data_out <= 8'he6;
         4077: data_out <= 8'h04;
         4078: data_out <= 8'h4f;
         4079: data_out <= 8'h58;
         4080: data_out <= 8'hcb;
         4081: data_out <= 8'h05;
         4082: data_out <= 8'hbd;
         4083: data_out <= 8'h03;
         4084: data_out <= 8'h12;
         4085: data_out <= 8'h9c;
         4086: data_out <= 8'ha3;
         4087: data_out <= 8'h27;
         4088: data_out <= 8'hdf;
         4089: data_out <= 8'h8d;
         4090: data_out <= 8'h08;
         4091: data_out <= 8'h20;
         4092: data_out <= 8'hf8;
         4093: data_out <= 8'ha6;
         4094: data_out <= 8'h01;
         4095: data_out <= 8'h08;
         4096: data_out <= 8'h08;
         4097: data_out <= 8'h2a;
         4098: data_out <= 8'h22;
         4099: data_out <= 8'he6;
         4100: data_out <= 8'h00;
         4101: data_out <= 8'h27;
         4102: data_out <= 8'h1e;
         4103: data_out <= 8'ha6;
         4104: data_out <= 8'h02;
         4105: data_out <= 8'h91;
         4106: data_out <= 8'h84;
         4107: data_out <= 8'h22;
         4108: data_out <= 8'h18;
         4109: data_out <= 8'he6;
         4110: data_out <= 8'h03;
         4111: data_out <= 8'h25;
         4112: data_out <= 8'h04;
         4113: data_out <= 8'hd1;
         4114: data_out <= 8'h85;
         4115: data_out <= 8'h24;
         4116: data_out <= 8'h10;
         4117: data_out <= 8'h91;
         4118: data_out <= 8'ha9;
         4119: data_out <= 8'h25;
         4120: data_out <= 8'h0c;
         4121: data_out <= 8'h22;
         4122: data_out <= 8'h04;
         4123: data_out <= 8'hd1;
         4124: data_out <= 8'haa;
         4125: data_out <= 8'h23;
         4126: data_out <= 8'h06;
         4127: data_out <= 8'hdf;
         4128: data_out <= 8'hab;
         4129: data_out <= 8'h97;
         4130: data_out <= 8'ha9;
         4131: data_out <= 8'hd7;
         4132: data_out <= 8'haa;
         4133: data_out <= 8'h08;
         4134: data_out <= 8'h08;
         4135: data_out <= 8'h08;
         4136: data_out <= 8'h08;
         4137: data_out <= 8'h39;
         4138: data_out <= 8'hde;
         4139: data_out <= 8'hab;
         4140: data_out <= 8'h27;
         4141: data_out <= 8'hfb;
         4142: data_out <= 8'h4f;
         4143: data_out <= 8'he6;
         4144: data_out <= 8'h00;
         4145: data_out <= 8'h5a;
         4146: data_out <= 8'hdb;
         4147: data_out <= 8'haa;
         4148: data_out <= 8'h99;
         4149: data_out <= 8'ha9;
         4150: data_out <= 8'h97;
         4151: data_out <= 8'ha5;
         4152: data_out <= 8'hd7;
         4153: data_out <= 8'ha6;
         4154: data_out <= 8'hde;
         4155: data_out <= 8'h84;
         4156: data_out <= 8'hdf;
         4157: data_out <= 8'ha3;
         4158: data_out <= 8'hbd;
         4159: data_out <= 8'h02;
         4160: data_out <= 8'hde;
         4161: data_out <= 8'hde;
         4162: data_out <= 8'hab;
         4163: data_out <= 8'h96;
         4164: data_out <= 8'ha7;
         4165: data_out <= 8'hd6;
         4166: data_out <= 8'ha8;
         4167: data_out <= 8'ha7;
         4168: data_out <= 8'h02;
         4169: data_out <= 8'he7;
         4170: data_out <= 8'h03;
         4171: data_out <= 8'hde;
         4172: data_out <= 8'ha7;
         4173: data_out <= 8'h09;
         4174: data_out <= 8'h7e;
         4175: data_out <= 8'h0f;
         4176: data_out <= 8'hb4;
         4177: data_out <= 8'h96;
         4178: data_out <= 8'hb2;
         4179: data_out <= 8'h36;
         4180: data_out <= 8'h96;
         4181: data_out <= 8'hb1;
         4182: data_out <= 8'h36;
         4183: data_out <= 8'hbd;
         4184: data_out <= 8'h0a;
         4185: data_out <= 8'hf9;
         4186: data_out <= 8'hbd;
         4187: data_out <= 8'h0a;
         4188: data_out <= 8'h1c;
         4189: data_out <= 8'h32;
         4190: data_out <= 8'h97;
         4191: data_out <= 8'hbb;
         4192: data_out <= 8'h32;
         4193: data_out <= 8'h97;
         4194: data_out <= 8'hbc;
         4195: data_out <= 8'hde;
         4196: data_out <= 8'hbb;
         4197: data_out <= 8'he6;
         4198: data_out <= 8'h00;
         4199: data_out <= 8'hde;
         4200: data_out <= 8'hb1;
         4201: data_out <= 8'heb;
         4202: data_out <= 8'h00;
         4203: data_out <= 8'h24;
         4204: data_out <= 8'h05;
         4205: data_out <= 8'hc6;
         4206: data_out <= 8'h1c;
         4207: data_out <= 8'h7e;
         4208: data_out <= 8'h03;
         4209: data_out <= 8'h21;
         4210: data_out <= 8'hbd;
         4211: data_out <= 8'h0f;
         4212: data_out <= 8'h2d;
         4213: data_out <= 8'hde;
         4214: data_out <= 8'hbb;
         4215: data_out <= 8'he6;
         4216: data_out <= 8'h00;
         4217: data_out <= 8'h8d;
         4218: data_out <= 8'h10;
         4219: data_out <= 8'hde;
         4220: data_out <= 8'had;
         4221: data_out <= 8'h8d;
         4222: data_out <= 8'h2c;
         4223: data_out <= 8'h8d;
         4224: data_out <= 8'h0c;
         4225: data_out <= 8'hde;
         4226: data_out <= 8'hbb;
         4227: data_out <= 8'h8d;
         4228: data_out <= 8'h26;
         4229: data_out <= 8'hbd;
         4230: data_out <= 8'h0f;
         4231: data_out <= 8'h66;
         4232: data_out <= 8'h7e;
         4233: data_out <= 8'h0a;
         4234: data_out <= 8'h3b;
         4235: data_out <= 8'hee;
         4236: data_out <= 8'h02;
         4237: data_out <= 8'h07;
         4238: data_out <= 8'h36;
         4239: data_out <= 8'h9f;
         4240: data_out <= 8'h78;
         4241: data_out <= 8'h0f;
         4242: data_out <= 8'h35;
         4243: data_out <= 8'hde;
         4244: data_out <= 8'h86;
         4245: data_out <= 8'h5c;
         4246: data_out <= 8'h20;
         4247: data_out <= 8'h04;
         4248: data_out <= 8'h32;
         4249: data_out <= 8'ha7;
         4250: data_out <= 8'h00;
         4251: data_out <= 8'h08;
         4252: data_out <= 8'h5a;
         4253: data_out <= 8'h26;
         4254: data_out <= 8'hf9;
         4255: data_out <= 8'hdf;
         4256: data_out <= 8'h86;
         4257: data_out <= 8'h9e;
         4258: data_out <= 8'h78;
         4259: data_out <= 8'h32;
         4260: data_out <= 8'h06;
         4261: data_out <= 8'h39;
         4262: data_out <= 8'hbd;
         4263: data_out <= 8'h0a;
         4264: data_out <= 8'h1c;
         4265: data_out <= 8'hde;
         4266: data_out <= 8'hb1;
         4267: data_out <= 8'he6;
         4268: data_out <= 8'h00;
         4269: data_out <= 8'h8d;
         4270: data_out <= 8'h18;
         4271: data_out <= 8'h26;
         4272: data_out <= 8'h13;
         4273: data_out <= 8'hee;
         4274: data_out <= 8'h06;
         4275: data_out <= 8'h09;
         4276: data_out <= 8'h9c;
         4277: data_out <= 8'h84;
         4278: data_out <= 8'h26;
         4279: data_out <= 8'h0a;
         4280: data_out <= 8'h37;
         4281: data_out <= 8'hdb;
         4282: data_out <= 8'h85;
         4283: data_out <= 8'h99;
         4284: data_out <= 8'h84;
         4285: data_out <= 8'h97;
         4286: data_out <= 8'h84;
         4287: data_out <= 8'hd7;
         4288: data_out <= 8'h85;
         4289: data_out <= 8'h33;
         4290: data_out <= 8'h08;
         4291: data_out <= 8'h39;
         4292: data_out <= 8'hee;
         4293: data_out <= 8'h02;
         4294: data_out <= 8'h39;
         4295: data_out <= 8'h9c;
         4296: data_out <= 8'h63;
         4297: data_out <= 8'h26;
         4298: data_out <= 8'h09;
         4299: data_out <= 8'hdf;
         4300: data_out <= 8'h61;
         4301: data_out <= 8'h09;
         4302: data_out <= 8'h09;
         4303: data_out <= 8'h09;
         4304: data_out <= 8'h09;
         4305: data_out <= 8'hdf;
         4306: data_out <= 8'h63;
         4307: data_out <= 8'h4f;
         4308: data_out <= 8'h39;
         4309: data_out <= 8'h8d;
         4310: data_out <= 8'h03;
         4311: data_out <= 8'h7e;
         4312: data_out <= 8'h0e;
         4313: data_out <= 8'h6e;
         4314: data_out <= 8'h8d;
         4315: data_out <= 8'hca;
         4316: data_out <= 8'h7f;
         4317: data_out <= 8'h00;
         4318: data_out <= 8'h5c;
         4319: data_out <= 8'h5d;
         4320: data_out <= 8'h39;
         4321: data_out <= 8'hbd;
         4322: data_out <= 8'h11;
         4323: data_out <= 8'h6d;
         4324: data_out <= 8'hc6;
         4325: data_out <= 8'h01;
         4326: data_out <= 8'hbd;
         4327: data_out <= 8'h0f;
         4328: data_out <= 8'h84;
         4329: data_out <= 8'h96;
         4330: data_out <= 8'hb2;
         4331: data_out <= 8'hbd;
         4332: data_out <= 8'h0f;
         4333: data_out <= 8'h31;
         4334: data_out <= 8'ha7;
         4335: data_out <= 8'h00;
         4336: data_out <= 8'h31;
         4337: data_out <= 8'h31;
         4338: data_out <= 8'h7e;
         4339: data_out <= 8'h0f;
         4340: data_out <= 8'h66;
         4341: data_out <= 8'h8d;
         4342: data_out <= 8'h02;
         4343: data_out <= 8'h20;
         4344: data_out <= 8'hde;
         4345: data_out <= 8'h8d;
         4346: data_out <= 8'hdf;
         4347: data_out <= 8'h27;
         4348: data_out <= 8'h67;
         4349: data_out <= 8'he6;
         4350: data_out <= 8'h00;
         4351: data_out <= 8'h39;
         4352: data_out <= 8'h8d;
         4353: data_out <= 8'h45;
         4354: data_out <= 8'h4f;
         4355: data_out <= 8'he1;
         4356: data_out <= 8'h00;
         4357: data_out <= 8'h23;
         4358: data_out <= 8'h03;
         4359: data_out <= 8'he6;
         4360: data_out <= 8'h00;
         4361: data_out <= 8'h4f;
         4362: data_out <= 8'h37;
         4363: data_out <= 8'h36;
         4364: data_out <= 8'hbd;
         4365: data_out <= 8'h0f;
         4366: data_out <= 8'h2f;
         4367: data_out <= 8'hde;
         4368: data_out <= 8'had;
         4369: data_out <= 8'h8d;
         4370: data_out <= 8'h98;
         4371: data_out <= 8'h33;
         4372: data_out <= 8'hbd;
         4373: data_out <= 8'h03;
         4374: data_out <= 8'h11;
         4375: data_out <= 8'h33;
         4376: data_out <= 8'hbd;
         4377: data_out <= 8'h10;
         4378: data_out <= 8'h8d;
         4379: data_out <= 8'h20;
         4380: data_out <= 8'hd5;
         4381: data_out <= 8'h8d;
         4382: data_out <= 8'h28;
         4383: data_out <= 8'ha6;
         4384: data_out <= 8'h00;
         4385: data_out <= 8'h10;
         4386: data_out <= 8'h20;
         4387: data_out <= 8'hdf;
         4388: data_out <= 8'hc6;
         4389: data_out <= 8'hff;
         4390: data_out <= 8'hd7;
         4391: data_out <= 8'hb2;
         4392: data_out <= 8'h8d;
         4393: data_out <= 8'h4c;
         4394: data_out <= 8'h81;
         4395: data_out <= 8'h29;
         4396: data_out <= 8'h27;
         4397: data_out <= 8'h05;
         4398: data_out <= 8'hbd;
         4399: data_out <= 8'h0b;
         4400: data_out <= 8'h4b;
         4401: data_out <= 8'h8d;
         4402: data_out <= 8'h37;
         4403: data_out <= 8'h8d;
         4404: data_out <= 8'h12;
         4405: data_out <= 8'h5f;
         4406: data_out <= 8'h4a;
         4407: data_out <= 8'ha1;
         4408: data_out <= 8'h00;
         4409: data_out <= 8'h24;
         4410: data_out <= 8'hcf;
         4411: data_out <= 8'h16;
         4412: data_out <= 8'he0;
         4413: data_out <= 8'h00;
         4414: data_out <= 8'h50;
         4415: data_out <= 8'hd1;
         4416: data_out <= 8'hb2;
         4417: data_out <= 8'h23;
         4418: data_out <= 8'hc7;
         4419: data_out <= 8'hd6;
         4420: data_out <= 8'hb2;
         4421: data_out <= 8'h20;
         4422: data_out <= 8'hc3;
         4423: data_out <= 8'hbd;
         4424: data_out <= 8'h0b;
         4425: data_out <= 8'h45;
         4426: data_out <= 8'h33;
         4427: data_out <= 8'hd7;
         4428: data_out <= 8'h78;
         4429: data_out <= 8'h33;
         4430: data_out <= 8'hd7;
         4431: data_out <= 8'h79;
         4432: data_out <= 8'h31;
         4433: data_out <= 8'h31;
         4434: data_out <= 8'h32;
         4435: data_out <= 8'h33;
         4436: data_out <= 8'hd7;
         4437: data_out <= 8'had;
         4438: data_out <= 8'h33;
         4439: data_out <= 8'hd7;
         4440: data_out <= 8'hae;
         4441: data_out <= 8'hde;
         4442: data_out <= 8'had;
         4443: data_out <= 8'hd6;
         4444: data_out <= 8'h79;
         4445: data_out <= 8'h37;
         4446: data_out <= 8'hd6;
         4447: data_out <= 8'h78;
         4448: data_out <= 8'h37;
         4449: data_out <= 8'h16;
         4450: data_out <= 8'h26;
         4451: data_out <= 8'h3b;
         4452: data_out <= 8'h7e;
         4453: data_out <= 8'h0d;
         4454: data_out <= 8'h71;
         4455: data_out <= 8'hbd;
         4456: data_out <= 8'h00;
         4457: data_out <= 8'hbf;
         4458: data_out <= 8'hbd;
         4459: data_out <= 8'h0a;
         4460: data_out <= 8'h19;
         4461: data_out <= 8'hbd;
         4462: data_out <= 8'h0c;
         4463: data_out <= 8'hea;
         4464: data_out <= 8'h96;
         4465: data_out <= 8'hb1;
         4466: data_out <= 8'h26;
         4467: data_out <= 8'hf0;
         4468: data_out <= 8'hd6;
         4469: data_out <= 8'hb2;
         4470: data_out <= 8'h7e;
         4471: data_out <= 8'h00;
         4472: data_out <= 8'hc7;
         4473: data_out <= 8'hbd;
         4474: data_out <= 8'h10;
         4475: data_out <= 8'hda;
         4476: data_out <= 8'h26;
         4477: data_out <= 8'h03;
         4478: data_out <= 8'h7e;
         4479: data_out <= 8'h13;
         4480: data_out <= 8'h85;
         4481: data_out <= 8'hbd;
         4482: data_out <= 8'h03;
         4483: data_out <= 8'h11;
         4484: data_out <= 8'ha6;
         4485: data_out <= 8'h00;
         4486: data_out <= 8'h36;
         4487: data_out <= 8'h6f;
         4488: data_out <= 8'h00;
         4489: data_out <= 8'hde;
         4490: data_out <= 8'hc8;
         4491: data_out <= 8'hdf;
         4492: data_out <= 8'hbd;
         4493: data_out <= 8'hde;
         4494: data_out <= 8'h71;
         4495: data_out <= 8'hdf;
         4496: data_out <= 8'hc8;
         4497: data_out <= 8'h8d;
         4498: data_out <= 8'he3;
         4499: data_out <= 8'hbd;
         4500: data_out <= 8'h16;
         4501: data_out <= 8'h7c;
         4502: data_out <= 8'h32;
         4503: data_out <= 8'hde;
         4504: data_out <= 8'h73;
         4505: data_out <= 8'ha7;
         4506: data_out <= 8'h00;
         4507: data_out <= 8'hde;
         4508: data_out <= 8'hbd;
         4509: data_out <= 8'hdf;
         4510: data_out <= 8'hc8;
         4511: data_out <= 8'h39;
         4512: data_out <= 8'hbd;
         4513: data_out <= 8'h0a;
         4514: data_out <= 8'h19;
         4515: data_out <= 8'h8d;
         4516: data_out <= 8'h07;
         4517: data_out <= 8'hdf;
         4518: data_out <= 8'h8e;
         4519: data_out <= 8'hbd;
         4520: data_out <= 8'h0b;
         4521: data_out <= 8'h4b;
         4522: data_out <= 8'h20;
         4523: data_out <= 8'hbe;
         4524: data_out <= 8'h96;
         4525: data_out <= 8'hb3;
         4526: data_out <= 8'h2b;
         4527: data_out <= 8'hb4;
         4528: data_out <= 8'h96;
         4529: data_out <= 8'haf;
         4530: data_out <= 8'h81;
         4531: data_out <= 8'h90;
         4532: data_out <= 8'h22;
         4533: data_out <= 8'hae;
         4534: data_out <= 8'hbd;
         4535: data_out <= 8'h16;
         4536: data_out <= 8'h30;
         4537: data_out <= 8'hde;
         4538: data_out <= 8'hb1;
         4539: data_out <= 8'h39;
         4540: data_out <= 8'h8d;
         4541: data_out <= 8'hee;
         4542: data_out <= 8'he6;
         4543: data_out <= 8'h00;
         4544: data_out <= 8'h7e;
         4545: data_out <= 8'h0e;
         4546: data_out <= 8'h6e;
         4547: data_out <= 8'h8d;
         4548: data_out <= 8'hdb;
         4549: data_out <= 8'hde;
         4550: data_out <= 8'h8e;
         4551: data_out <= 8'he7;
         4552: data_out <= 8'h00;
         4553: data_out <= 8'h39;
         4554: data_out <= 8'h8d;
         4555: data_out <= 8'hd4;
         4556: data_out <= 8'hd7;
         4557: data_out <= 8'h9e;
         4558: data_out <= 8'h5f;
         4559: data_out <= 8'hbd;
         4560: data_out <= 8'h00;
         4561: data_out <= 8'hc7;
         4562: data_out <= 8'h27;
         4563: data_out <= 8'h02;
         4564: data_out <= 8'h8d;
         4565: data_out <= 8'hd1;
         4566: data_out <= 8'hd7;
         4567: data_out <= 8'h9f;
         4568: data_out <= 8'hde;
         4569: data_out <= 8'h8e;
         4570: data_out <= 8'ha6;
         4571: data_out <= 8'h00;
         4572: data_out <= 8'h98;
         4573: data_out <= 8'h9f;
         4574: data_out <= 8'h94;
         4575: data_out <= 8'h9e;
         4576: data_out <= 8'h27;
         4577: data_out <= 8'hf8;
         4578: data_out <= 8'h39;
         4579: data_out <= 8'h81;
         4580: data_out <= 8'ha5;
         4581: data_out <= 8'h26;
         4582: data_out <= 8'h03;
         4583: data_out <= 8'h7e;
         4584: data_out <= 8'h12;
         4585: data_out <= 8'ha5;
         4586: data_out <= 8'hbd;
         4587: data_out <= 8'h0a;
         4588: data_out <= 8'h27;
         4589: data_out <= 8'hbd;
         4590: data_out <= 8'h10;
         4591: data_out <= 8'hf9;
         4592: data_out <= 8'h86;
         4593: data_out <= 8'hd3;
         4594: data_out <= 8'hbd;
         4595: data_out <= 8'h12;
         4596: data_out <= 8'h78;
         4597: data_out <= 8'h8d;
         4598: data_out <= 8'h7f;
         4599: data_out <= 8'h17;
         4600: data_out <= 8'h8d;
         4601: data_out <= 8'h7e;
         4602: data_out <= 8'hde;
         4603: data_out <= 8'h7a;
         4604: data_out <= 8'ha6;
         4605: data_out <= 8'h00;
         4606: data_out <= 8'h08;
         4607: data_out <= 8'h8d;
         4608: data_out <= 8'h77;
         4609: data_out <= 8'h9c;
         4610: data_out <= 8'h7c;
         4611: data_out <= 8'h26;
         4612: data_out <= 8'hf7;
         4613: data_out <= 8'h39;
         4614: data_out <= 8'h81;
         4615: data_out <= 8'ha5;
         4616: data_out <= 8'h26;
         4617: data_out <= 8'h03;
         4618: data_out <= 8'h7e;
         4619: data_out <= 8'h12;
         4620: data_out <= 8'ha8;
         4621: data_out <= 8'h7f;
         4622: data_out <= 8'h00;
         4623: data_out <= 8'hb0;
         4624: data_out <= 8'h81;
         4625: data_out <= 8'h97;
         4626: data_out <= 8'h26;
         4627: data_out <= 8'h08;
         4628: data_out <= 8'h7a;
         4629: data_out <= 8'h00;
         4630: data_out <= 8'hb0;
         4631: data_out <= 8'hde;
         4632: data_out <= 8'hc8;
         4633: data_out <= 8'h08;
         4634: data_out <= 8'hdf;
         4635: data_out <= 8'hc8;
         4636: data_out <= 8'hbd;
         4637: data_out <= 8'h0a;
         4638: data_out <= 8'h27;
         4639: data_out <= 8'hbd;
         4640: data_out <= 8'h10;
         4641: data_out <= 8'hf9;
         4642: data_out <= 8'h96;
         4643: data_out <= 8'hb0;
         4644: data_out <= 8'h26;
         4645: data_out <= 8'h03;
         4646: data_out <= 8'hbd;
         4647: data_out <= 8'h04;
         4648: data_out <= 8'hf2;
         4649: data_out <= 8'h37;
         4650: data_out <= 8'hc6;
         4651: data_out <= 8'h03;
         4652: data_out <= 8'h8d;
         4653: data_out <= 8'h55;
         4654: data_out <= 8'h81;
         4655: data_out <= 8'hd3;
         4656: data_out <= 8'h26;
         4657: data_out <= 8'hf8;
         4658: data_out <= 8'h5a;
         4659: data_out <= 8'h26;
         4660: data_out <= 8'hf7;
         4661: data_out <= 8'h8d;
         4662: data_out <= 8'h4c;
         4663: data_out <= 8'h33;
         4664: data_out <= 8'h11;
         4665: data_out <= 8'h26;
         4666: data_out <= 8'hee;
         4667: data_out <= 8'hde;
         4668: data_out <= 8'h7a;
         4669: data_out <= 8'h09;
         4670: data_out <= 8'h20;
         4671: data_out <= 8'h1b;
         4672: data_out <= 8'h8d;
         4673: data_out <= 8'h41;
         4674: data_out <= 8'ha7;
         4675: data_out <= 8'h00;
         4676: data_out <= 8'h8d;
         4677: data_out <= 8'h48;
         4678: data_out <= 8'ha7;
         4679: data_out <= 8'h00;
         4680: data_out <= 8'h8d;
         4681: data_out <= 8'h44;
         4682: data_out <= 8'ha7;
         4683: data_out <= 8'h00;
         4684: data_out <= 8'hdf;
         4685: data_out <= 8'hb1;
         4686: data_out <= 8'h96;
         4687: data_out <= 8'hb1;
         4688: data_out <= 8'hd6;
         4689: data_out <= 8'hb2;
         4690: data_out <= 8'hbd;
         4691: data_out <= 8'h02;
         4692: data_out <= 8'hfe;
         4693: data_out <= 8'h8d;
         4694: data_out <= 8'h37;
         4695: data_out <= 8'ha7;
         4696: data_out <= 8'h00;
         4697: data_out <= 8'h26;
         4698: data_out <= 8'hf1;
         4699: data_out <= 8'h8d;
         4700: data_out <= 8'h26;
         4701: data_out <= 8'ha7;
         4702: data_out <= 8'h00;
         4703: data_out <= 8'h26;
         4704: data_out <= 8'hdf;
         4705: data_out <= 8'h8d;
         4706: data_out <= 8'h20;
         4707: data_out <= 8'ha7;
         4708: data_out <= 8'h00;
         4709: data_out <= 8'h26;
         4710: data_out <= 8'hdd;
         4711: data_out <= 8'h08;
         4712: data_out <= 8'hdf;
         4713: data_out <= 8'h7c;
         4714: data_out <= 8'hce;
         4715: data_out <= 8'h02;
         4716: data_out <= 8'ha5;
         4717: data_out <= 8'hbd;
         4718: data_out <= 8'h08;
         4719: data_out <= 8'h87;
         4720: data_out <= 8'hbd;
         4721: data_out <= 8'h03;
         4722: data_out <= 8'hd0;
         4723: data_out <= 8'h7e;
         4724: data_out <= 8'h03;
         4725: data_out <= 8'h53;
         4726: data_out <= 8'h8d;
         4727: data_out <= 8'h00;
         4728: data_out <= 8'h36;
         4729: data_out <= 8'hb6;
         4730: data_out <= 8'hf0;
         4731: data_out <= 8'h10;
         4732: data_out <= 8'h2b;
         4733: data_out <= 8'hfb;
         4734: data_out <= 8'h32;
         4735: data_out <= 8'hb7;
         4736: data_out <= 8'hf0;
         4737: data_out <= 8'h11;
         4738: data_out <= 8'h39;
         4739: data_out <= 8'hb6;
         4740: data_out <= 8'hf0;
         4741: data_out <= 8'h10;
         4742: data_out <= 8'h46;
         4743: data_out <= 8'h25;
         4744: data_out <= 8'hfa;
         4745: data_out <= 8'h08;
         4746: data_out <= 8'hb6;
         4747: data_out <= 8'hf0;
         4748: data_out <= 8'h11;
         4749: data_out <= 8'h39;
         4750: data_out <= 8'h8d;
         4751: data_out <= 8'hf3;
         4752: data_out <= 8'h36;
         4753: data_out <= 8'ha0;
         4754: data_out <= 8'h00;
         4755: data_out <= 8'h94;
         4756: data_out <= 8'hb0;
         4757: data_out <= 8'h32;
         4758: data_out <= 8'h26;
         4759: data_out <= 8'h01;
         4760: data_out <= 8'h39;
         4761: data_out <= 8'hce;
         4762: data_out <= 8'h12;
         4763: data_out <= 8'hfd;
         4764: data_out <= 8'hbd;
         4765: data_out <= 8'h08;
         4766: data_out <= 8'h87;
         4767: data_out <= 8'hbd;
         4768: data_out <= 8'h05;
         4769: data_out <= 8'h0e;
         4770: data_out <= 8'h7e;
         4771: data_out <= 8'h03;
         4772: data_out <= 8'h4a;
         4773: data_out <= 8'hc6;
         4774: data_out <= 8'hff;
         4775: data_out <= 8'h86;
         4776: data_out <= 8'h5f;
         4777: data_out <= 8'h37;
         4778: data_out <= 8'hbd;
         4779: data_out <= 8'h00;
         4780: data_out <= 8'hbf;
         4781: data_out <= 8'hc6;
         4782: data_out <= 8'h01;
         4783: data_out <= 8'hd7;
         4784: data_out <= 8'h5e;
         4785: data_out <= 8'h7e;
         4786: data_out <= 8'h0c;
         4787: data_out <= 8'h37;
         4788: data_out <= 8'hbd;
         4789: data_out <= 8'h0a;
         4790: data_out <= 8'h1d;
         4791: data_out <= 8'ha6;
         4792: data_out <= 8'h02;
         4793: data_out <= 8'he6;
         4794: data_out <= 8'h03;
         4795: data_out <= 8'hbd;
         4796: data_out <= 8'h03;
         4797: data_out <= 8'h12;
         4798: data_out <= 8'hde;
         4799: data_out <= 8'h71;
         4800: data_out <= 8'he6;
         4801: data_out <= 8'h04;
         4802: data_out <= 8'h58;
         4803: data_out <= 8'hcb;
         4804: data_out <= 8'h05;
         4805: data_out <= 8'hdb;
         4806: data_out <= 8'h72;
         4807: data_out <= 8'h4f;
         4808: data_out <= 8'h99;
         4809: data_out <= 8'h71;
         4810: data_out <= 8'h97;
         4811: data_out <= 8'h71;
         4812: data_out <= 8'hd7;
         4813: data_out <= 8'h72;
         4814: data_out <= 8'h32;
         4815: data_out <= 8'h97;
         4816: data_out <= 8'hb1;
         4817: data_out <= 8'h26;
         4818: data_out <= 8'h0d;
         4819: data_out <= 8'hc6;
         4820: data_out <= 8'h04;
         4821: data_out <= 8'h8d;
         4822: data_out <= 8'hac;
         4823: data_out <= 8'h81;
         4824: data_out <= 8'hd2;
         4825: data_out <= 8'h26;
         4826: data_out <= 8'hf8;
         4827: data_out <= 8'h5a;
         4828: data_out <= 8'h26;
         4829: data_out <= 8'hf7;
         4830: data_out <= 8'h20;
         4831: data_out <= 8'h06;
         4832: data_out <= 8'h86;
         4833: data_out <= 8'hd2;
         4834: data_out <= 8'h8d;
         4835: data_out <= 8'h92;
         4836: data_out <= 8'h8d;
         4837: data_out <= 8'h90;
         4838: data_out <= 8'hde;
         4839: data_out <= 8'h71;
         4840: data_out <= 8'h9c;
         4841: data_out <= 8'h73;
         4842: data_out <= 8'h27;
         4843: data_out <= 8'ha1;
         4844: data_out <= 8'ha6;
         4845: data_out <= 8'h00;
         4846: data_out <= 8'hd6;
         4847: data_out <= 8'hb1;
         4848: data_out <= 8'h27;
         4849: data_out <= 8'h04;
         4850: data_out <= 8'h8d;
         4851: data_out <= 8'h84;
         4852: data_out <= 8'h20;
         4853: data_out <= 8'h05;
         4854: data_out <= 8'h8d;
         4855: data_out <= 8'h8b;
         4856: data_out <= 8'h09;
         4857: data_out <= 8'ha7;
         4858: data_out <= 8'h00;
         4859: data_out <= 8'h08;
         4860: data_out <= 8'h20;
         4861: data_out <= 8'hea;
         4862: data_out <= 8'h4e;
         4863: data_out <= 8'h4f;
         4864: data_out <= 8'h20;
         4865: data_out <= 8'h47;
         4866: data_out <= 8'h4f;
         4867: data_out <= 8'h4f;
         4868: data_out <= 8'h44;
         4869: data_out <= 8'h09;
         4870: data_out <= 8'h89;
         4871: data_out <= 8'h0d;
         4872: data_out <= 8'h0a;
         4873: data_out <= 8'h00;
         4874: data_out <= 8'hce;
         4875: data_out <= 8'h18;
         4876: data_out <= 8'h3c;
         4877: data_out <= 8'h20;
         4878: data_out <= 8'h0b;
         4879: data_out <= 8'hbd;
         4880: data_out <= 8'h14;
         4881: data_out <= 8'hab;
         4882: data_out <= 8'h73;
         4883: data_out <= 8'h00;
         4884: data_out <= 8'hb3;
         4885: data_out <= 8'h73;
         4886: data_out <= 8'h00;
         4887: data_out <= 8'hbb;
         4888: data_out <= 8'h20;
         4889: data_out <= 8'h03;
         4890: data_out <= 8'hbd;
         4891: data_out <= 8'h14;
         4892: data_out <= 8'hab;
         4893: data_out <= 8'h5d;
         4894: data_out <= 8'h26;
         4895: data_out <= 8'h03;
         4896: data_out <= 8'h7e;
         4897: data_out <= 8'h15;
         4898: data_out <= 8'hbf;
         4899: data_out <= 8'hce;
         4900: data_out <= 8'h00;
         4901: data_out <= 8'hb6;
         4902: data_out <= 8'h16;
         4903: data_out <= 8'h27;
         4904: data_out <= 8'h61;
         4905: data_out <= 8'hd0;
         4906: data_out <= 8'haf;
         4907: data_out <= 8'h27;
         4908: data_out <= 8'h5e;
         4909: data_out <= 8'h2b;
         4910: data_out <= 8'h0a;
         4911: data_out <= 8'h97;
         4912: data_out <= 8'haf;
         4913: data_out <= 8'h96;
         4914: data_out <= 8'hba;
         4915: data_out <= 8'h97;
         4916: data_out <= 8'hb3;
         4917: data_out <= 8'hce;
         4918: data_out <= 8'h00;
         4919: data_out <= 8'haf;
         4920: data_out <= 8'h50;
         4921: data_out <= 8'hc1;
         4922: data_out <= 8'hf8;
         4923: data_out <= 8'h2f;
         4924: data_out <= 8'h4e;
         4925: data_out <= 8'h4f;
         4926: data_out <= 8'h64;
         4927: data_out <= 8'h01;
         4928: data_out <= 8'hbd;
         4929: data_out <= 8'h13;
         4930: data_out <= 8'hfe;
         4931: data_out <= 8'hd6;
         4932: data_out <= 8'hbb;
         4933: data_out <= 8'h2a;
         4934: data_out <= 8'h09;
         4935: data_out <= 8'h63;
         4936: data_out <= 8'h01;
         4937: data_out <= 8'h63;
         4938: data_out <= 8'h02;
         4939: data_out <= 8'h63;
         4940: data_out <= 8'h03;
         4941: data_out <= 8'h43;
         4942: data_out <= 8'h89;
         4943: data_out <= 8'h00;
         4944: data_out <= 8'h97;
         4945: data_out <= 8'hbc;
         4946: data_out <= 8'h96;
         4947: data_out <= 8'hb2;
         4948: data_out <= 8'h99;
         4949: data_out <= 8'hb9;
         4950: data_out <= 8'h97;
         4951: data_out <= 8'hb2;
         4952: data_out <= 8'h96;
         4953: data_out <= 8'hb1;
         4954: data_out <= 8'h99;
         4955: data_out <= 8'hb8;
         4956: data_out <= 8'h97;
         4957: data_out <= 8'hb1;
         4958: data_out <= 8'h96;
         4959: data_out <= 8'hb0;
         4960: data_out <= 8'h99;
         4961: data_out <= 8'hb7;
         4962: data_out <= 8'h97;
         4963: data_out <= 8'hb0;
         4964: data_out <= 8'h17;
         4965: data_out <= 8'h2a;
         4966: data_out <= 8'h40;
         4967: data_out <= 8'h25;
         4968: data_out <= 8'h02;
         4969: data_out <= 8'h8d;
         4970: data_out <= 8'h58;
         4971: data_out <= 8'h5f;
         4972: data_out <= 8'h96;
         4973: data_out <= 8'hb0;
         4974: data_out <= 8'h26;
         4975: data_out <= 8'h2d;
         4976: data_out <= 8'h96;
         4977: data_out <= 8'hb1;
         4978: data_out <= 8'h97;
         4979: data_out <= 8'hb0;
         4980: data_out <= 8'h96;
         4981: data_out <= 8'hb2;
         4982: data_out <= 8'h97;
         4983: data_out <= 8'hb1;
         4984: data_out <= 8'h96;
         4985: data_out <= 8'hbc;
         4986: data_out <= 8'h97;
         4987: data_out <= 8'hb2;
         4988: data_out <= 8'h7f;
         4989: data_out <= 8'h00;
         4990: data_out <= 8'hbc;
         4991: data_out <= 8'hcb;
         4992: data_out <= 8'h08;
         4993: data_out <= 8'hc1;
         4994: data_out <= 8'h20;
         4995: data_out <= 8'h2d;
         4996: data_out <= 8'he7;
         4997: data_out <= 8'h4f;
         4998: data_out <= 8'h97;
         4999: data_out <= 8'haf;
         5000: data_out <= 8'h97;
         5001: data_out <= 8'hb3;
         5002: data_out <= 8'h39;
         5003: data_out <= 8'h8d;
         5004: data_out <= 8'h65;
         5005: data_out <= 8'h0c;
         5006: data_out <= 8'h20;
         5007: data_out <= 8'hb3;
         5008: data_out <= 8'h5c;
         5009: data_out <= 8'h78;
         5010: data_out <= 8'h00;
         5011: data_out <= 8'hbc;
         5012: data_out <= 8'h79;
         5013: data_out <= 8'h00;
         5014: data_out <= 8'hb2;
         5015: data_out <= 8'h79;
         5016: data_out <= 8'h00;
         5017: data_out <= 8'hb1;
         5018: data_out <= 8'h79;
         5019: data_out <= 8'h00;
         5020: data_out <= 8'hb0;
         5021: data_out <= 8'h2a;
         5022: data_out <= 8'hf1;
         5023: data_out <= 8'h96;
         5024: data_out <= 8'haf;
         5025: data_out <= 8'h10;
         5026: data_out <= 8'h97;
         5027: data_out <= 8'haf;
         5028: data_out <= 8'h23;
         5029: data_out <= 8'hdf;
         5030: data_out <= 8'h8c;
         5031: data_out <= 8'h25;
         5032: data_out <= 8'h05;
         5033: data_out <= 8'h78;
         5034: data_out <= 8'h00;
         5035: data_out <= 8'hbc;
         5036: data_out <= 8'h20;
         5037: data_out <= 8'h0e;
         5038: data_out <= 8'h7c;
         5039: data_out <= 8'h00;
         5040: data_out <= 8'haf;
         5041: data_out <= 8'h27;
         5042: data_out <= 8'h27;
         5043: data_out <= 8'h76;
         5044: data_out <= 8'h00;
         5045: data_out <= 8'hb0;
         5046: data_out <= 8'h76;
         5047: data_out <= 8'h00;
         5048: data_out <= 8'hb1;
         5049: data_out <= 8'h76;
         5050: data_out <= 8'h00;
         5051: data_out <= 8'hb2;
         5052: data_out <= 8'h24;
         5053: data_out <= 8'h04;
         5054: data_out <= 8'h8d;
         5055: data_out <= 8'h0f;
         5056: data_out <= 8'h27;
         5057: data_out <= 8'hec;
         5058: data_out <= 8'h39;
         5059: data_out <= 8'h73;
         5060: data_out <= 8'h00;
         5061: data_out <= 8'hb3;
         5062: data_out <= 8'h73;
         5063: data_out <= 8'h00;
         5064: data_out <= 8'hb0;
         5065: data_out <= 8'h73;
         5066: data_out <= 8'h00;
         5067: data_out <= 8'hb1;
         5068: data_out <= 8'h73;
         5069: data_out <= 8'h00;
         5070: data_out <= 8'hb2;
         5071: data_out <= 8'hde;
         5072: data_out <= 8'hb1;
         5073: data_out <= 8'h08;
         5074: data_out <= 8'hdf;
         5075: data_out <= 8'hb1;
         5076: data_out <= 8'h26;
         5077: data_out <= 8'h03;
         5078: data_out <= 8'h7c;
         5079: data_out <= 8'h00;
         5080: data_out <= 8'hb0;
         5081: data_out <= 8'h39;
         5082: data_out <= 8'hc6;
         5083: data_out <= 8'h0a;
         5084: data_out <= 8'h7e;
         5085: data_out <= 8'h03;
         5086: data_out <= 8'h21;
         5087: data_out <= 8'hce;
         5088: data_out <= 8'h00;
         5089: data_out <= 8'h74;
         5090: data_out <= 8'ha6;
         5091: data_out <= 8'h03;
         5092: data_out <= 8'h97;
         5093: data_out <= 8'hbc;
         5094: data_out <= 8'ha6;
         5095: data_out <= 8'h02;
         5096: data_out <= 8'ha7;
         5097: data_out <= 8'h03;
         5098: data_out <= 8'ha6;
         5099: data_out <= 8'h01;
         5100: data_out <= 8'ha7;
         5101: data_out <= 8'h02;
         5102: data_out <= 8'h96;
         5103: data_out <= 8'hb5;
         5104: data_out <= 8'ha7;
         5105: data_out <= 8'h01;
         5106: data_out <= 8'hcb;
         5107: data_out <= 8'h08;
         5108: data_out <= 8'h2f;
         5109: data_out <= 8'hec;
         5110: data_out <= 8'h96;
         5111: data_out <= 8'hbc;
         5112: data_out <= 8'hc0;
         5113: data_out <= 8'h08;
         5114: data_out <= 8'h27;
         5115: data_out <= 8'h0a;
         5116: data_out <= 8'h67;
         5117: data_out <= 8'h01;
         5118: data_out <= 8'h66;
         5119: data_out <= 8'h02;
         5120: data_out <= 8'h66;
         5121: data_out <= 8'h03;
         5122: data_out <= 8'h46;
         5123: data_out <= 8'h5c;
         5124: data_out <= 8'h26;
         5125: data_out <= 8'hf6;
         5126: data_out <= 8'h39;
         5127: data_out <= 8'h81;
         5128: data_out <= 8'h00;
         5129: data_out <= 8'h00;
         5130: data_out <= 8'h00;
         5131: data_out <= 8'h02;
         5132: data_out <= 8'h80;
         5133: data_out <= 8'h19;
         5134: data_out <= 8'h56;
         5135: data_out <= 8'haa;
         5136: data_out <= 8'h80;
         5137: data_out <= 8'h76;
         5138: data_out <= 8'h22;
         5139: data_out <= 8'hf1;
         5140: data_out <= 8'h82;
         5141: data_out <= 8'h38;
         5142: data_out <= 8'haa;
         5143: data_out <= 8'h45;
         5144: data_out <= 8'h80;
         5145: data_out <= 8'h35;
         5146: data_out <= 8'h04;
         5147: data_out <= 8'hf3;
         5148: data_out <= 8'h81;
         5149: data_out <= 8'h35;
         5150: data_out <= 8'h04;
         5151: data_out <= 8'hf3;
         5152: data_out <= 8'h80;
         5153: data_out <= 8'h80;
         5154: data_out <= 8'h00;
         5155: data_out <= 8'h00;
         5156: data_out <= 8'h80;
         5157: data_out <= 8'h31;
         5158: data_out <= 8'h72;
         5159: data_out <= 8'h18;
         5160: data_out <= 8'hbd;
         5161: data_out <= 8'h15;
         5162: data_out <= 8'hd9;
         5163: data_out <= 8'h2e;
         5164: data_out <= 8'h03;
         5165: data_out <= 8'h7e;
         5166: data_out <= 8'h0d;
         5167: data_out <= 8'h71;
         5168: data_out <= 8'hce;
         5169: data_out <= 8'h14;
         5170: data_out <= 8'h18;
         5171: data_out <= 8'h96;
         5172: data_out <= 8'haf;
         5173: data_out <= 8'h80;
         5174: data_out <= 8'h80;
         5175: data_out <= 8'h36;
         5176: data_out <= 8'h86;
         5177: data_out <= 8'h80;
         5178: data_out <= 8'h97;
         5179: data_out <= 8'haf;
         5180: data_out <= 8'hbd;
         5181: data_out <= 8'h13;
         5182: data_out <= 8'h1a;
         5183: data_out <= 8'hce;
         5184: data_out <= 8'h14;
         5185: data_out <= 8'h1c;
         5186: data_out <= 8'hbd;
         5187: data_out <= 8'h15;
         5188: data_out <= 8'h12;
         5189: data_out <= 8'hce;
         5190: data_out <= 8'h14;
         5191: data_out <= 8'h07;
         5192: data_out <= 8'hbd;
         5193: data_out <= 8'h13;
         5194: data_out <= 8'h0f;
         5195: data_out <= 8'hce;
         5196: data_out <= 8'h14;
         5197: data_out <= 8'h0b;
         5198: data_out <= 8'hbd;
         5199: data_out <= 8'h18;
         5200: data_out <= 8'hf7;
         5201: data_out <= 8'hce;
         5202: data_out <= 8'h14;
         5203: data_out <= 8'h20;
         5204: data_out <= 8'hbd;
         5205: data_out <= 8'h13;
         5206: data_out <= 8'h1a;
         5207: data_out <= 8'h33;
         5208: data_out <= 8'hbd;
         5209: data_out <= 8'h17;
         5210: data_out <= 8'h07;
         5211: data_out <= 8'hce;
         5212: data_out <= 8'h14;
         5213: data_out <= 8'h24;
         5214: data_out <= 8'h8d;
         5215: data_out <= 8'h4b;
         5216: data_out <= 8'h27;
         5217: data_out <= 8'h48;
         5218: data_out <= 8'h8d;
         5219: data_out <= 8'h63;
         5220: data_out <= 8'h86;
         5221: data_out <= 8'h00;
         5222: data_out <= 8'h97;
         5223: data_out <= 8'h75;
         5224: data_out <= 8'h97;
         5225: data_out <= 8'h76;
         5226: data_out <= 8'h97;
         5227: data_out <= 8'h77;
         5228: data_out <= 8'hd6;
         5229: data_out <= 8'hb2;
         5230: data_out <= 8'h8d;
         5231: data_out <= 8'h0e;
         5232: data_out <= 8'hd6;
         5233: data_out <= 8'hb1;
         5234: data_out <= 8'h8d;
         5235: data_out <= 8'h0a;
         5236: data_out <= 8'hd6;
         5237: data_out <= 8'hb0;
         5238: data_out <= 8'h8d;
         5239: data_out <= 8'h0b;
         5240: data_out <= 8'hbd;
         5241: data_out <= 8'h15;
         5242: data_out <= 8'h85;
         5243: data_out <= 8'h7e;
         5244: data_out <= 8'h13;
         5245: data_out <= 8'h6b;
         5246: data_out <= 8'h26;
         5247: data_out <= 8'h03;
         5248: data_out <= 8'h7e;
         5249: data_out <= 8'h13;
         5250: data_out <= 8'hdf;
         5251: data_out <= 8'h0d;
         5252: data_out <= 8'h96;
         5253: data_out <= 8'h75;
         5254: data_out <= 8'h56;
         5255: data_out <= 8'h27;
         5256: data_out <= 8'h21;
         5257: data_out <= 8'h24;
         5258: data_out <= 8'h10;
         5259: data_out <= 8'h96;
         5260: data_out <= 8'h77;
         5261: data_out <= 8'h9b;
         5262: data_out <= 8'hb9;
         5263: data_out <= 8'h97;
         5264: data_out <= 8'h77;
         5265: data_out <= 8'h96;
         5266: data_out <= 8'h76;
         5267: data_out <= 8'h99;
         5268: data_out <= 8'hb8;
         5269: data_out <= 8'h97;
         5270: data_out <= 8'h76;
         5271: data_out <= 8'h96;
         5272: data_out <= 8'h75;
         5273: data_out <= 8'h99;
         5274: data_out <= 8'hb7;
         5275: data_out <= 8'h46;
         5276: data_out <= 8'h97;
         5277: data_out <= 8'h75;
         5278: data_out <= 8'h76;
         5279: data_out <= 8'h00;
         5280: data_out <= 8'h76;
         5281: data_out <= 8'h76;
         5282: data_out <= 8'h00;
         5283: data_out <= 8'h77;
         5284: data_out <= 8'h76;
         5285: data_out <= 8'h00;
         5286: data_out <= 8'hbc;
         5287: data_out <= 8'h0c;
         5288: data_out <= 8'h20;
         5289: data_out <= 8'hda;
         5290: data_out <= 8'h39;
         5291: data_out <= 8'ha6;
         5292: data_out <= 8'h01;
         5293: data_out <= 8'h97;
         5294: data_out <= 8'hba;
         5295: data_out <= 8'h16;
         5296: data_out <= 8'h8a;
         5297: data_out <= 8'h80;
         5298: data_out <= 8'h97;
         5299: data_out <= 8'hb7;
         5300: data_out <= 8'hd8;
         5301: data_out <= 8'hb3;
         5302: data_out <= 8'hd7;
         5303: data_out <= 8'hbb;
         5304: data_out <= 8'ha6;
         5305: data_out <= 8'h02;
         5306: data_out <= 8'h97;
         5307: data_out <= 8'hb8;
         5308: data_out <= 8'ha6;
         5309: data_out <= 8'h03;
         5310: data_out <= 8'h97;
         5311: data_out <= 8'hb9;
         5312: data_out <= 8'ha6;
         5313: data_out <= 8'h00;
         5314: data_out <= 8'h97;
         5315: data_out <= 8'hb6;
         5316: data_out <= 8'hd6;
         5317: data_out <= 8'haf;
         5318: data_out <= 8'h39;
         5319: data_out <= 8'h4d;
         5320: data_out <= 8'h27;
         5321: data_out <= 8'h19;
         5322: data_out <= 8'h9b;
         5323: data_out <= 8'haf;
         5324: data_out <= 8'h46;
         5325: data_out <= 8'h49;
         5326: data_out <= 8'h28;
         5327: data_out <= 8'h13;
         5328: data_out <= 8'h8b;
         5329: data_out <= 8'h80;
         5330: data_out <= 8'h97;
         5331: data_out <= 8'haf;
         5332: data_out <= 8'h26;
         5333: data_out <= 8'h03;
         5334: data_out <= 8'h7e;
         5335: data_out <= 8'h13;
         5336: data_out <= 8'h88;
         5337: data_out <= 8'h96;
         5338: data_out <= 8'hbb;
         5339: data_out <= 8'h97;
         5340: data_out <= 8'hb3;
         5341: data_out <= 8'h39;
         5342: data_out <= 8'h96;
         5343: data_out <= 8'hb3;
         5344: data_out <= 8'h43;
         5345: data_out <= 8'h20;
         5346: data_out <= 8'h02;
         5347: data_out <= 8'h32;
         5348: data_out <= 8'h32;
         5349: data_out <= 8'h2b;
         5350: data_out <= 8'h03;
         5351: data_out <= 8'h7e;
         5352: data_out <= 8'h13;
         5353: data_out <= 8'h85;
         5354: data_out <= 8'h7e;
         5355: data_out <= 8'h13;
         5356: data_out <= 8'hda;
         5357: data_out <= 8'hbd;
         5358: data_out <= 8'h15;
         5359: data_out <= 8'hcc;
         5360: data_out <= 8'h27;
         5361: data_out <= 8'h0f;
         5362: data_out <= 8'h8b;
         5363: data_out <= 8'h02;
         5364: data_out <= 8'h25;
         5365: data_out <= 8'hf4;
         5366: data_out <= 8'h7f;
         5367: data_out <= 8'h00;
         5368: data_out <= 8'hbb;
         5369: data_out <= 8'hbd;
         5370: data_out <= 8'h13;
         5371: data_out <= 8'h26;
         5372: data_out <= 8'h7c;
         5373: data_out <= 8'h00;
         5374: data_out <= 8'haf;
         5375: data_out <= 8'h27;
         5376: data_out <= 8'he9;
         5377: data_out <= 8'h39;
         5378: data_out <= 8'h84;
         5379: data_out <= 8'h20;
         5380: data_out <= 8'h00;
         5381: data_out <= 8'h00;
         5382: data_out <= 8'hbd;
         5383: data_out <= 8'h15;
         5384: data_out <= 8'hcc;
         5385: data_out <= 8'hce;
         5386: data_out <= 8'h15;
         5387: data_out <= 8'h02;
         5388: data_out <= 8'h5f;
         5389: data_out <= 8'hd7;
         5390: data_out <= 8'hbb;
         5391: data_out <= 8'h8d;
         5392: data_out <= 8'h7d;
         5393: data_out <= 8'h8c;
         5394: data_out <= 8'h8d;
         5395: data_out <= 8'h97;
         5396: data_out <= 8'h27;
         5397: data_out <= 8'h6a;
         5398: data_out <= 8'h70;
         5399: data_out <= 8'h00;
         5400: data_out <= 8'haf;
         5401: data_out <= 8'h8d;
         5402: data_out <= 8'hac;
         5403: data_out <= 8'h7c;
         5404: data_out <= 8'h00;
         5405: data_out <= 8'haf;
         5406: data_out <= 8'h27;
         5407: data_out <= 8'hca;
         5408: data_out <= 8'hce;
         5409: data_out <= 8'h00;
         5410: data_out <= 8'h75;
         5411: data_out <= 8'hc6;
         5412: data_out <= 8'h03;
         5413: data_out <= 8'hd7;
         5414: data_out <= 8'h5a;
         5415: data_out <= 8'hc6;
         5416: data_out <= 8'h01;
         5417: data_out <= 8'h96;
         5418: data_out <= 8'hb0;
         5419: data_out <= 8'h91;
         5420: data_out <= 8'hb7;
         5421: data_out <= 8'h26;
         5422: data_out <= 8'h0d;
         5423: data_out <= 8'h96;
         5424: data_out <= 8'hb1;
         5425: data_out <= 8'h91;
         5426: data_out <= 8'hb8;
         5427: data_out <= 8'h26;
         5428: data_out <= 8'h07;
         5429: data_out <= 8'h96;
         5430: data_out <= 8'hb2;
         5431: data_out <= 8'h91;
         5432: data_out <= 8'hb9;
         5433: data_out <= 8'h26;
         5434: data_out <= 8'h01;
         5435: data_out <= 8'h0d;
         5436: data_out <= 8'h07;
         5437: data_out <= 8'h59;
         5438: data_out <= 8'h24;
         5439: data_out <= 8'h0c;
         5440: data_out <= 8'he7;
         5441: data_out <= 8'h00;
         5442: data_out <= 8'h08;
         5443: data_out <= 8'h7a;
         5444: data_out <= 8'h00;
         5445: data_out <= 8'h5a;
         5446: data_out <= 8'h2b;
         5447: data_out <= 8'h2e;
         5448: data_out <= 8'h27;
         5449: data_out <= 8'h28;
         5450: data_out <= 8'hc6;
         5451: data_out <= 8'h01;
         5452: data_out <= 8'h06;
         5453: data_out <= 8'h25;
         5454: data_out <= 8'h0f;
         5455: data_out <= 8'h78;
         5456: data_out <= 8'h00;
         5457: data_out <= 8'hb9;
         5458: data_out <= 8'h79;
         5459: data_out <= 8'h00;
         5460: data_out <= 8'hb8;
         5461: data_out <= 8'h79;
         5462: data_out <= 8'h00;
         5463: data_out <= 8'hb7;
         5464: data_out <= 8'h25;
         5465: data_out <= 8'he2;
         5466: data_out <= 8'h2b;
         5467: data_out <= 8'hcd;
         5468: data_out <= 8'h20;
         5469: data_out <= 8'hde;
         5470: data_out <= 8'h96;
         5471: data_out <= 8'hb9;
         5472: data_out <= 8'h90;
         5473: data_out <= 8'hb2;
         5474: data_out <= 8'h97;
         5475: data_out <= 8'hb9;
         5476: data_out <= 8'h96;
         5477: data_out <= 8'hb8;
         5478: data_out <= 8'h92;
         5479: data_out <= 8'hb1;
         5480: data_out <= 8'h97;
         5481: data_out <= 8'hb8;
         5482: data_out <= 8'h96;
         5483: data_out <= 8'hb7;
         5484: data_out <= 8'h92;
         5485: data_out <= 8'hb0;
         5486: data_out <= 8'h97;
         5487: data_out <= 8'hb7;
         5488: data_out <= 8'h20;
         5489: data_out <= 8'hdd;
         5490: data_out <= 8'hc6;
         5491: data_out <= 8'h40;
         5492: data_out <= 8'h20;
         5493: data_out <= 8'hd6;
         5494: data_out <= 8'h56;
         5495: data_out <= 8'h56;
         5496: data_out <= 8'h56;
         5497: data_out <= 8'hd7;
         5498: data_out <= 8'hbc;
         5499: data_out <= 8'h8d;
         5500: data_out <= 8'h08;
         5501: data_out <= 8'h7e;
         5502: data_out <= 8'h13;
         5503: data_out <= 8'h6b;
         5504: data_out <= 8'hc6;
         5505: data_out <= 8'h14;
         5506: data_out <= 8'h7e;
         5507: data_out <= 8'h03;
         5508: data_out <= 8'h21;
         5509: data_out <= 8'hde;
         5510: data_out <= 8'h75;
         5511: data_out <= 8'hdf;
         5512: data_out <= 8'hb0;
         5513: data_out <= 8'h96;
         5514: data_out <= 8'h77;
         5515: data_out <= 8'h97;
         5516: data_out <= 8'hb2;
         5517: data_out <= 8'h39;
         5518: data_out <= 8'he6;
         5519: data_out <= 8'h01;
         5520: data_out <= 8'hd7;
         5521: data_out <= 8'hb3;
         5522: data_out <= 8'hca;
         5523: data_out <= 8'h80;
         5524: data_out <= 8'hd7;
         5525: data_out <= 8'hb0;
         5526: data_out <= 8'he6;
         5527: data_out <= 8'h00;
         5528: data_out <= 8'hee;
         5529: data_out <= 8'h02;
         5530: data_out <= 8'hdf;
         5531: data_out <= 8'hb1;
         5532: data_out <= 8'hd7;
         5533: data_out <= 8'haf;
         5534: data_out <= 8'h39;
         5535: data_out <= 8'hce;
         5536: data_out <= 8'h00;
         5537: data_out <= 8'ha7;
         5538: data_out <= 8'h20;
         5539: data_out <= 8'h06;
         5540: data_out <= 8'hce;
         5541: data_out <= 8'h00;
         5542: data_out <= 8'ha3;
         5543: data_out <= 8'h8c;
         5544: data_out <= 8'hde;
         5545: data_out <= 8'h9e;
         5546: data_out <= 8'h96;
         5547: data_out <= 8'haf;
         5548: data_out <= 8'ha7;
         5549: data_out <= 8'h00;
         5550: data_out <= 8'h96;
         5551: data_out <= 8'hb3;
         5552: data_out <= 8'h8a;
         5553: data_out <= 8'h7f;
         5554: data_out <= 8'h94;
         5555: data_out <= 8'hb0;
         5556: data_out <= 8'ha7;
         5557: data_out <= 8'h01;
         5558: data_out <= 8'h96;
         5559: data_out <= 8'hb1;
         5560: data_out <= 8'ha7;
         5561: data_out <= 8'h02;
         5562: data_out <= 8'h96;
         5563: data_out <= 8'hb2;
         5564: data_out <= 8'ha7;
         5565: data_out <= 8'h03;
         5566: data_out <= 8'h39;
         5567: data_out <= 8'h96;
         5568: data_out <= 8'hba;
         5569: data_out <= 8'h97;
         5570: data_out <= 8'hb3;
         5571: data_out <= 8'hde;
         5572: data_out <= 8'hb6;
         5573: data_out <= 8'hdf;
         5574: data_out <= 8'haf;
         5575: data_out <= 8'hde;
         5576: data_out <= 8'hb8;
         5577: data_out <= 8'hdf;
         5578: data_out <= 8'hb1;
         5579: data_out <= 8'h39;
         5580: data_out <= 8'hde;
         5581: data_out <= 8'hb0;
         5582: data_out <= 8'hdf;
         5583: data_out <= 8'hb7;
         5584: data_out <= 8'hde;
         5585: data_out <= 8'hb2;
         5586: data_out <= 8'hdf;
         5587: data_out <= 8'hb9;
         5588: data_out <= 8'h96;
         5589: data_out <= 8'haf;
         5590: data_out <= 8'h97;
         5591: data_out <= 8'hb6;
         5592: data_out <= 8'h39;
         5593: data_out <= 8'hd6;
         5594: data_out <= 8'haf;
         5595: data_out <= 8'h27;
         5596: data_out <= 8'h08;
         5597: data_out <= 8'hd6;
         5598: data_out <= 8'hb3;
         5599: data_out <= 8'h59;
         5600: data_out <= 8'hc6;
         5601: data_out <= 8'hff;
         5602: data_out <= 8'h25;
         5603: data_out <= 8'h01;
         5604: data_out <= 8'h50;
         5605: data_out <= 8'h39;
         5606: data_out <= 8'h8d;
         5607: data_out <= 8'hf1;
         5608: data_out <= 8'hd7;
         5609: data_out <= 8'hb0;
         5610: data_out <= 8'h7f;
         5611: data_out <= 8'h00;
         5612: data_out <= 8'hb1;
         5613: data_out <= 8'hc6;
         5614: data_out <= 8'h88;
         5615: data_out <= 8'h96;
         5616: data_out <= 8'hb0;
         5617: data_out <= 8'h80;
         5618: data_out <= 8'h80;
         5619: data_out <= 8'hd7;
         5620: data_out <= 8'haf;
         5621: data_out <= 8'h86;
         5622: data_out <= 8'h00;
         5623: data_out <= 8'h97;
         5624: data_out <= 8'hb2;
         5625: data_out <= 8'h97;
         5626: data_out <= 8'hbc;
         5627: data_out <= 8'h97;
         5628: data_out <= 8'hb3;
         5629: data_out <= 8'h7e;
         5630: data_out <= 8'h13;
         5631: data_out <= 8'h67;
         5632: data_out <= 8'h7f;
         5633: data_out <= 8'h00;
         5634: data_out <= 8'hb3;
         5635: data_out <= 8'h39;
         5636: data_out <= 8'he6;
         5637: data_out <= 8'h00;
         5638: data_out <= 8'h27;
         5639: data_out <= 8'hd1;
         5640: data_out <= 8'he6;
         5641: data_out <= 8'h01;
         5642: data_out <= 8'hd8;
         5643: data_out <= 8'hb3;
         5644: data_out <= 8'h2b;
         5645: data_out <= 8'hcf;
         5646: data_out <= 8'hd6;
         5647: data_out <= 8'haf;
         5648: data_out <= 8'he1;
         5649: data_out <= 8'h00;
         5650: data_out <= 8'h26;
         5651: data_out <= 8'h17;
         5652: data_out <= 8'he6;
         5653: data_out <= 8'h01;
         5654: data_out <= 8'hca;
         5655: data_out <= 8'h7f;
         5656: data_out <= 8'hd4;
         5657: data_out <= 8'hb0;
         5658: data_out <= 8'he1;
         5659: data_out <= 8'h01;
         5660: data_out <= 8'h26;
         5661: data_out <= 8'h0d;
         5662: data_out <= 8'hd6;
         5663: data_out <= 8'hb1;
         5664: data_out <= 8'he1;
         5665: data_out <= 8'h02;
         5666: data_out <= 8'h26;
         5667: data_out <= 8'h07;
         5668: data_out <= 8'hd6;
         5669: data_out <= 8'hb2;
         5670: data_out <= 8'he0;
         5671: data_out <= 8'h03;
         5672: data_out <= 8'h26;
         5673: data_out <= 8'h01;
         5674: data_out <= 8'h39;
         5675: data_out <= 8'h56;
         5676: data_out <= 8'hd8;
         5677: data_out <= 8'hb3;
         5678: data_out <= 8'h20;
         5679: data_out <= 8'haf;
         5680: data_out <= 8'hd6;
         5681: data_out <= 8'haf;
         5682: data_out <= 8'h27;
         5683: data_out <= 8'h41;
         5684: data_out <= 8'hc0;
         5685: data_out <= 8'h98;
         5686: data_out <= 8'h96;
         5687: data_out <= 8'hb3;
         5688: data_out <= 8'h2a;
         5689: data_out <= 8'h06;
         5690: data_out <= 8'h73;
         5691: data_out <= 8'h00;
         5692: data_out <= 8'hb5;
         5693: data_out <= 8'hbd;
         5694: data_out <= 8'h13;
         5695: data_out <= 8'hc6;
         5696: data_out <= 8'hce;
         5697: data_out <= 8'h00;
         5698: data_out <= 8'haf;
         5699: data_out <= 8'hc1;
         5700: data_out <= 8'hf8;
         5701: data_out <= 8'h2e;
         5702: data_out <= 8'h07;
         5703: data_out <= 8'hbd;
         5704: data_out <= 8'h13;
         5705: data_out <= 8'hf2;
         5706: data_out <= 8'h7f;
         5707: data_out <= 8'h00;
         5708: data_out <= 8'hb5;
         5709: data_out <= 8'h39;
         5710: data_out <= 8'h7f;
         5711: data_out <= 8'h00;
         5712: data_out <= 8'hb5;
         5713: data_out <= 8'h96;
         5714: data_out <= 8'hb3;
         5715: data_out <= 8'h49;
         5716: data_out <= 8'h76;
         5717: data_out <= 8'h00;
         5718: data_out <= 8'hb0;
         5719: data_out <= 8'h7e;
         5720: data_out <= 8'h13;
         5721: data_out <= 8'hfe;
         5722: data_out <= 8'hd6;
         5723: data_out <= 8'haf;
         5724: data_out <= 8'hc1;
         5725: data_out <= 8'h98;
         5726: data_out <= 8'h24;
         5727: data_out <= 8'h1b;
         5728: data_out <= 8'h8d;
         5729: data_out <= 8'hce;
         5730: data_out <= 8'hd7;
         5731: data_out <= 8'hbc;
         5732: data_out <= 8'h96;
         5733: data_out <= 8'hb3;
         5734: data_out <= 8'hd7;
         5735: data_out <= 8'hb3;
         5736: data_out <= 8'h80;
         5737: data_out <= 8'h80;
         5738: data_out <= 8'h86;
         5739: data_out <= 8'h98;
         5740: data_out <= 8'h97;
         5741: data_out <= 8'haf;
         5742: data_out <= 8'h96;
         5743: data_out <= 8'hb2;
         5744: data_out <= 8'h97;
         5745: data_out <= 8'h58;
         5746: data_out <= 8'h7e;
         5747: data_out <= 8'h13;
         5748: data_out <= 8'h67;
         5749: data_out <= 8'hd7;
         5750: data_out <= 8'hb0;
         5751: data_out <= 8'hd7;
         5752: data_out <= 8'hb1;
         5753: data_out <= 8'hd7;
         5754: data_out <= 8'hb2;
         5755: data_out <= 8'h39;
         5756: data_out <= 8'hce;
         5757: data_out <= 8'h00;
         5758: data_out <= 8'h00;
         5759: data_out <= 8'hdf;
         5760: data_out <= 8'hb3;
         5761: data_out <= 8'hdf;
         5762: data_out <= 8'haf;
         5763: data_out <= 8'hdf;
         5764: data_out <= 8'hb1;
         5765: data_out <= 8'hdf;
         5766: data_out <= 8'ha9;
         5767: data_out <= 8'hdf;
         5768: data_out <= 8'ha7;
         5769: data_out <= 8'h25;
         5770: data_out <= 8'h6b;
         5771: data_out <= 8'h81;
         5772: data_out <= 8'h2d;
         5773: data_out <= 8'h26;
         5774: data_out <= 8'h05;
         5775: data_out <= 8'h73;
         5776: data_out <= 8'h00;
         5777: data_out <= 8'hb4;
         5778: data_out <= 8'h20;
         5779: data_out <= 8'h04;
         5780: data_out <= 8'h81;
         5781: data_out <= 8'h2b;
         5782: data_out <= 8'h26;
         5783: data_out <= 8'h05;
         5784: data_out <= 8'hbd;
         5785: data_out <= 8'h00;
         5786: data_out <= 8'hbf;
         5787: data_out <= 8'h25;
         5788: data_out <= 8'h59;
         5789: data_out <= 8'h81;
         5790: data_out <= 8'h2e;
         5791: data_out <= 8'h27;
         5792: data_out <= 8'h2d;
         5793: data_out <= 8'h81;
         5794: data_out <= 8'h45;
         5795: data_out <= 8'h26;
         5796: data_out <= 8'h2e;
         5797: data_out <= 8'hbd;
         5798: data_out <= 8'h00;
         5799: data_out <= 8'hbf;
         5800: data_out <= 8'h25;
         5801: data_out <= 8'h69;
         5802: data_out <= 8'h81;
         5803: data_out <= 8'ha4;
         5804: data_out <= 8'h27;
         5805: data_out <= 8'h0e;
         5806: data_out <= 8'h81;
         5807: data_out <= 8'h2d;
         5808: data_out <= 8'h27;
         5809: data_out <= 8'h0a;
         5810: data_out <= 8'h81;
         5811: data_out <= 8'ha3;
         5812: data_out <= 8'h27;
         5813: data_out <= 8'h09;
         5814: data_out <= 8'h81;
         5815: data_out <= 8'h2b;
         5816: data_out <= 8'h27;
         5817: data_out <= 8'h05;
         5818: data_out <= 8'h20;
         5819: data_out <= 8'h08;
         5820: data_out <= 8'h73;
         5821: data_out <= 8'h00;
         5822: data_out <= 8'haa;
         5823: data_out <= 8'hbd;
         5824: data_out <= 8'h00;
         5825: data_out <= 8'hbf;
         5826: data_out <= 8'h25;
         5827: data_out <= 8'h4f;
         5828: data_out <= 8'h7d;
         5829: data_out <= 8'h00;
         5830: data_out <= 8'haa;
         5831: data_out <= 8'h27;
         5832: data_out <= 8'h0a;
         5833: data_out <= 8'h70;
         5834: data_out <= 8'h00;
         5835: data_out <= 8'ha9;
         5836: data_out <= 8'h20;
         5837: data_out <= 8'h05;
         5838: data_out <= 8'h73;
         5839: data_out <= 8'h00;
         5840: data_out <= 8'ha8;
         5841: data_out <= 8'h26;
         5842: data_out <= 8'hc5;
         5843: data_out <= 8'h96;
         5844: data_out <= 8'ha9;
         5845: data_out <= 8'h90;
         5846: data_out <= 8'ha7;
         5847: data_out <= 8'h97;
         5848: data_out <= 8'ha9;
         5849: data_out <= 8'h27;
         5850: data_out <= 8'h14;
         5851: data_out <= 8'h2a;
         5852: data_out <= 8'h0a;
         5853: data_out <= 8'hbd;
         5854: data_out <= 8'h15;
         5855: data_out <= 8'h06;
         5856: data_out <= 8'h7c;
         5857: data_out <= 8'h00;
         5858: data_out <= 8'ha9;
         5859: data_out <= 8'h26;
         5860: data_out <= 8'hf8;
         5861: data_out <= 8'h20;
         5862: data_out <= 8'h08;
         5863: data_out <= 8'hbd;
         5864: data_out <= 8'h14;
         5865: data_out <= 8'hed;
         5866: data_out <= 8'h7a;
         5867: data_out <= 8'h00;
         5868: data_out <= 8'ha9;
         5869: data_out <= 8'h26;
         5870: data_out <= 8'hf8;
         5871: data_out <= 8'h96;
         5872: data_out <= 8'hb4;
         5873: data_out <= 8'h2a;
         5874: data_out <= 8'h88;
         5875: data_out <= 8'h7e;
         5876: data_out <= 8'h18;
         5877: data_out <= 8'h91;
         5878: data_out <= 8'hd6;
         5879: data_out <= 8'ha7;
         5880: data_out <= 8'hd0;
         5881: data_out <= 8'ha8;
         5882: data_out <= 8'hd7;
         5883: data_out <= 8'ha7;
         5884: data_out <= 8'h36;
         5885: data_out <= 8'hbd;
         5886: data_out <= 8'h14;
         5887: data_out <= 8'hed;
         5888: data_out <= 8'h33;
         5889: data_out <= 8'hc0;
         5890: data_out <= 8'h30;
         5891: data_out <= 8'h8d;
         5892: data_out <= 8'h02;
         5893: data_out <= 8'h20;
         5894: data_out <= 8'h91;
         5895: data_out <= 8'hbd;
         5896: data_out <= 8'h15;
         5897: data_out <= 8'ha4;
         5898: data_out <= 8'hbd;
         5899: data_out <= 8'h15;
         5900: data_out <= 8'he8;
         5901: data_out <= 8'hce;
         5902: data_out <= 8'h00;
         5903: data_out <= 8'ha3;
         5904: data_out <= 8'h7e;
         5905: data_out <= 8'h13;
         5906: data_out <= 8'h1a;
         5907: data_out <= 8'hd6;
         5908: data_out <= 8'ha9;
         5909: data_out <= 8'h58;
         5910: data_out <= 8'h58;
         5911: data_out <= 8'hdb;
         5912: data_out <= 8'ha9;
         5913: data_out <= 8'h58;
         5914: data_out <= 8'h80;
         5915: data_out <= 8'h30;
         5916: data_out <= 8'h1b;
         5917: data_out <= 8'h97;
         5918: data_out <= 8'ha9;
         5919: data_out <= 8'h20;
         5920: data_out <= 8'h9e;
         5921: data_out <= 8'h91;
         5922: data_out <= 8'h43;
         5923: data_out <= 8'h4f;
         5924: data_out <= 8'hf8;
         5925: data_out <= 8'h94;
         5926: data_out <= 8'h74;
         5927: data_out <= 8'h23;
         5928: data_out <= 8'hf7;
         5929: data_out <= 8'h94;
         5930: data_out <= 8'h74;
         5931: data_out <= 8'h24;
         5932: data_out <= 8'h00;
         5933: data_out <= 8'hce;
         5934: data_out <= 8'h02;
         5935: data_out <= 8'ha0;
         5936: data_out <= 8'h8d;
         5937: data_out <= 8'h10;
         5938: data_out <= 8'h96;
         5939: data_out <= 8'h8a;
         5940: data_out <= 8'hd6;
         5941: data_out <= 8'h8b;
         5942: data_out <= 8'h97;
         5943: data_out <= 8'hb0;
         5944: data_out <= 8'hd7;
         5945: data_out <= 8'hb1;
         5946: data_out <= 8'hc6;
         5947: data_out <= 8'h90;
         5948: data_out <= 8'h0d;
         5949: data_out <= 8'hbd;
         5950: data_out <= 8'h15;
         5951: data_out <= 8'hf3;
         5952: data_out <= 8'h8d;
         5953: data_out <= 8'h03;
         5954: data_out <= 8'h7e;
         5955: data_out <= 8'h08;
         5956: data_out <= 8'h87;
         5957: data_out <= 8'hce;
         5958: data_out <= 8'h01;
         5959: data_out <= 8'h00;
         5960: data_out <= 8'h86;
         5961: data_out <= 8'h20;
         5962: data_out <= 8'hd6;
         5963: data_out <= 8'hb3;
         5964: data_out <= 8'h2a;
         5965: data_out <= 8'h02;
         5966: data_out <= 8'h86;
         5967: data_out <= 8'h2d;
         5968: data_out <= 8'ha7;
         5969: data_out <= 8'h00;
         5970: data_out <= 8'h97;
         5971: data_out <= 8'hb3;
         5972: data_out <= 8'hdf;
         5973: data_out <= 8'hbd;
         5974: data_out <= 8'h08;
         5975: data_out <= 8'h86;
         5976: data_out <= 8'h30;
         5977: data_out <= 8'hd6;
         5978: data_out <= 8'haf;
         5979: data_out <= 8'h26;
         5980: data_out <= 8'h03;
         5981: data_out <= 8'h7e;
         5982: data_out <= 8'h18;
         5983: data_out <= 8'h34;
         5984: data_out <= 8'h4f;
         5985: data_out <= 8'hc1;
         5986: data_out <= 8'h80;
         5987: data_out <= 8'h22;
         5988: data_out <= 8'h08;
         5989: data_out <= 8'hce;
         5990: data_out <= 8'h17;
         5991: data_out <= 8'h29;
         5992: data_out <= 8'hbd;
         5993: data_out <= 8'h14;
         5994: data_out <= 8'h5e;
         5995: data_out <= 8'h86;
         5996: data_out <= 8'hfa;
         5997: data_out <= 8'h97;
         5998: data_out <= 8'ha7;
         5999: data_out <= 8'hce;
         6000: data_out <= 8'h17;
         6001: data_out <= 8'h25;
         6002: data_out <= 8'hbd;
         6003: data_out <= 8'h16;
         6004: data_out <= 8'h0e;
         6005: data_out <= 8'h2e;
         6006: data_out <= 8'h10;
         6007: data_out <= 8'hce;
         6008: data_out <= 8'h17;
         6009: data_out <= 8'h21;
         6010: data_out <= 8'hbd;
         6011: data_out <= 8'h16;
         6012: data_out <= 8'h0e;
         6013: data_out <= 8'h2e;
         6014: data_out <= 8'h10;
         6015: data_out <= 8'hbd;
         6016: data_out <= 8'h14;
         6017: data_out <= 8'hed;
         6018: data_out <= 8'h7a;
         6019: data_out <= 8'h00;
         6020: data_out <= 8'ha7;
         6021: data_out <= 8'h20;
         6022: data_out <= 8'hf0;
         6023: data_out <= 8'hbd;
         6024: data_out <= 8'h15;
         6025: data_out <= 8'h06;
         6026: data_out <= 8'h7c;
         6027: data_out <= 8'h00;
         6028: data_out <= 8'ha7;
         6029: data_out <= 8'h20;
         6030: data_out <= 8'he0;
         6031: data_out <= 8'hbd;
         6032: data_out <= 8'h13;
         6033: data_out <= 8'h0a;
         6034: data_out <= 8'hbd;
         6035: data_out <= 8'h16;
         6036: data_out <= 8'h30;
         6037: data_out <= 8'hc6;
         6038: data_out <= 8'h01;
         6039: data_out <= 8'h96;
         6040: data_out <= 8'ha7;
         6041: data_out <= 8'h8b;
         6042: data_out <= 8'h07;
         6043: data_out <= 8'h2b;
         6044: data_out <= 8'h08;
         6045: data_out <= 8'h81;
         6046: data_out <= 8'h08;
         6047: data_out <= 8'h24;
         6048: data_out <= 8'h04;
         6049: data_out <= 8'h4a;
         6050: data_out <= 8'h16;
         6051: data_out <= 8'h86;
         6052: data_out <= 8'h02;
         6053: data_out <= 8'h4a;
         6054: data_out <= 8'h4a;
         6055: data_out <= 8'h97;
         6056: data_out <= 8'ha9;
         6057: data_out <= 8'hd7;
         6058: data_out <= 8'ha7;
         6059: data_out <= 8'h2e;
         6060: data_out <= 8'h11;
         6061: data_out <= 8'hde;
         6062: data_out <= 8'hbd;
         6063: data_out <= 8'h86;
         6064: data_out <= 8'h2e;
         6065: data_out <= 8'h08;
         6066: data_out <= 8'ha7;
         6067: data_out <= 8'h00;
         6068: data_out <= 8'h5d;
         6069: data_out <= 8'h27;
         6070: data_out <= 8'h05;
         6071: data_out <= 8'h86;
         6072: data_out <= 8'h30;
         6073: data_out <= 8'h08;
         6074: data_out <= 8'ha7;
         6075: data_out <= 8'h00;
         6076: data_out <= 8'hdf;
         6077: data_out <= 8'hbd;
         6078: data_out <= 8'hce;
         6079: data_out <= 8'h18;
         6080: data_out <= 8'h40;
         6081: data_out <= 8'hc6;
         6082: data_out <= 8'h80;
         6083: data_out <= 8'h96;
         6084: data_out <= 8'hb2;
         6085: data_out <= 8'hab;
         6086: data_out <= 8'h02;
         6087: data_out <= 8'h97;
         6088: data_out <= 8'hb2;
         6089: data_out <= 8'h96;
         6090: data_out <= 8'hb1;
         6091: data_out <= 8'ha9;
         6092: data_out <= 8'h01;
         6093: data_out <= 8'h97;
         6094: data_out <= 8'hb1;
         6095: data_out <= 8'h96;
         6096: data_out <= 8'hb0;
         6097: data_out <= 8'ha9;
         6098: data_out <= 8'h00;
         6099: data_out <= 8'h97;
         6100: data_out <= 8'hb0;
         6101: data_out <= 8'h5c;
         6102: data_out <= 8'h56;
         6103: data_out <= 8'h59;
         6104: data_out <= 8'h28;
         6105: data_out <= 8'he9;
         6106: data_out <= 8'h24;
         6107: data_out <= 8'h03;
         6108: data_out <= 8'hc0;
         6109: data_out <= 8'h0b;
         6110: data_out <= 8'h50;
         6111: data_out <= 8'hcb;
         6112: data_out <= 8'h2f;
         6113: data_out <= 8'h08;
         6114: data_out <= 8'h08;
         6115: data_out <= 8'h08;
         6116: data_out <= 8'hdf;
         6117: data_out <= 8'h9c;
         6118: data_out <= 8'hde;
         6119: data_out <= 8'hbd;
         6120: data_out <= 8'h08;
         6121: data_out <= 8'h17;
         6122: data_out <= 8'h84;
         6123: data_out <= 8'h7f;
         6124: data_out <= 8'ha7;
         6125: data_out <= 8'h00;
         6126: data_out <= 8'h7a;
         6127: data_out <= 8'h00;
         6128: data_out <= 8'ha7;
         6129: data_out <= 8'h26;
         6130: data_out <= 8'h05;
         6131: data_out <= 8'h86;
         6132: data_out <= 8'h2e;
         6133: data_out <= 8'h08;
         6134: data_out <= 8'ha7;
         6135: data_out <= 8'h00;
         6136: data_out <= 8'hdf;
         6137: data_out <= 8'hbd;
         6138: data_out <= 8'hde;
         6139: data_out <= 8'h9c;
         6140: data_out <= 8'h53;
         6141: data_out <= 8'hc4;
         6142: data_out <= 8'h80;
         6143: data_out <= 8'h8c;
         6144: data_out <= 8'h18;
         6145: data_out <= 8'h52;
         6146: data_out <= 8'h26;
         6147: data_out <= 8'hbf;
         6148: data_out <= 8'hde;
         6149: data_out <= 8'hbd;
         6150: data_out <= 8'ha6;
         6151: data_out <= 8'h00;
         6152: data_out <= 8'h09;
         6153: data_out <= 8'h81;
         6154: data_out <= 8'h30;
         6155: data_out <= 8'h27;
         6156: data_out <= 8'hf9;
         6157: data_out <= 8'h81;
         6158: data_out <= 8'h2e;
         6159: data_out <= 8'h27;
         6160: data_out <= 8'h01;
         6161: data_out <= 8'h08;
         6162: data_out <= 8'h86;
         6163: data_out <= 8'h2b;
         6164: data_out <= 8'hd6;
         6165: data_out <= 8'ha9;
         6166: data_out <= 8'h27;
         6167: data_out <= 8'h1e;
         6168: data_out <= 8'h2a;
         6169: data_out <= 8'h03;
         6170: data_out <= 8'h86;
         6171: data_out <= 8'h2d;
         6172: data_out <= 8'h50;
         6173: data_out <= 8'ha7;
         6174: data_out <= 8'h02;
         6175: data_out <= 8'h86;
         6176: data_out <= 8'h45;
         6177: data_out <= 8'ha7;
         6178: data_out <= 8'h01;
         6179: data_out <= 8'h86;
         6180: data_out <= 8'h2f;
         6181: data_out <= 8'h4c;
         6182: data_out <= 8'hc0;
         6183: data_out <= 8'h0a;
         6184: data_out <= 8'h24;
         6185: data_out <= 8'hfb;
         6186: data_out <= 8'hcb;
         6187: data_out <= 8'h3a;
         6188: data_out <= 8'ha7;
         6189: data_out <= 8'h03;
         6190: data_out <= 8'he7;
         6191: data_out <= 8'h04;
         6192: data_out <= 8'h6f;
         6193: data_out <= 8'h05;
         6194: data_out <= 8'h20;
         6195: data_out <= 8'h04;
         6196: data_out <= 8'ha7;
         6197: data_out <= 8'h00;
         6198: data_out <= 8'h6f;
         6199: data_out <= 8'h01;
         6200: data_out <= 8'hce;
         6201: data_out <= 8'h01;
         6202: data_out <= 8'h00;
         6203: data_out <= 8'h39;
         6204: data_out <= 8'h80;
         6205: data_out <= 8'h00;
         6206: data_out <= 8'h00;
         6207: data_out <= 8'h00;
         6208: data_out <= 8'hfe;
         6209: data_out <= 8'h79;
         6210: data_out <= 8'h60;
         6211: data_out <= 8'h00;
         6212: data_out <= 8'h27;
         6213: data_out <= 8'h10;
         6214: data_out <= 8'hff;
         6215: data_out <= 8'hfc;
         6216: data_out <= 8'h18;
         6217: data_out <= 8'h00;
         6218: data_out <= 8'h00;
         6219: data_out <= 8'h64;
         6220: data_out <= 8'hff;
         6221: data_out <= 8'hff;
         6222: data_out <= 8'hf6;
         6223: data_out <= 8'h00;
         6224: data_out <= 8'h00;
         6225: data_out <= 8'h01;
         6226: data_out <= 8'hbd;
         6227: data_out <= 8'h15;
         6228: data_out <= 8'hcc;
         6229: data_out <= 8'hce;
         6230: data_out <= 8'h18;
         6231: data_out <= 8'h3c;
         6232: data_out <= 8'hbd;
         6233: data_out <= 8'h15;
         6234: data_out <= 8'h8e;
         6235: data_out <= 8'h27;
         6236: data_out <= 8'h61;
         6237: data_out <= 8'h4d;
         6238: data_out <= 8'h26;
         6239: data_out <= 8'h03;
         6240: data_out <= 8'h7e;
         6241: data_out <= 8'h13;
         6242: data_out <= 8'h86;
         6243: data_out <= 8'hce;
         6244: data_out <= 8'h00;
         6245: data_out <= 8'hab;
         6246: data_out <= 8'hbd;
         6247: data_out <= 8'h15;
         6248: data_out <= 8'haa;
         6249: data_out <= 8'h5f;
         6250: data_out <= 8'h96;
         6251: data_out <= 8'hba;
         6252: data_out <= 8'h2a;
         6253: data_out <= 8'h10;
         6254: data_out <= 8'hbd;
         6255: data_out <= 8'h16;
         6256: data_out <= 8'h5a;
         6257: data_out <= 8'hce;
         6258: data_out <= 8'h00;
         6259: data_out <= 8'hab;
         6260: data_out <= 8'h96;
         6261: data_out <= 8'hba;
         6262: data_out <= 8'hbd;
         6263: data_out <= 8'h16;
         6264: data_out <= 8'h0e;
         6265: data_out <= 8'h26;
         6266: data_out <= 8'h03;
         6267: data_out <= 8'h43;
         6268: data_out <= 8'hd6;
         6269: data_out <= 8'h58;
         6270: data_out <= 8'hbd;
         6271: data_out <= 8'h15;
         6272: data_out <= 8'hc1;
         6273: data_out <= 8'h37;
         6274: data_out <= 8'hbd;
         6275: data_out <= 8'h14;
         6276: data_out <= 8'h28;
         6277: data_out <= 8'hce;
         6278: data_out <= 8'h00;
         6279: data_out <= 8'hab;
         6280: data_out <= 8'hbd;
         6281: data_out <= 8'h14;
         6282: data_out <= 8'h5e;
         6283: data_out <= 8'h8d;
         6284: data_out <= 8'h31;
         6285: data_out <= 8'h32;
         6286: data_out <= 8'h46;
         6287: data_out <= 8'h24;
         6288: data_out <= 8'haa;
         6289: data_out <= 8'h96;
         6290: data_out <= 8'haf;
         6291: data_out <= 8'h27;
         6292: data_out <= 8'h03;
         6293: data_out <= 8'h73;
         6294: data_out <= 8'h00;
         6295: data_out <= 8'hb3;
         6296: data_out <= 8'h39;
         6297: data_out <= 8'h81;
         6298: data_out <= 8'h38;
         6299: data_out <= 8'haa;
         6300: data_out <= 8'h3b;
         6301: data_out <= 8'h07;
         6302: data_out <= 8'h74;
         6303: data_out <= 8'h94;
         6304: data_out <= 8'h2e;
         6305: data_out <= 8'h40;
         6306: data_out <= 8'h77;
         6307: data_out <= 8'h2e;
         6308: data_out <= 8'h4f;
         6309: data_out <= 8'h70;
         6310: data_out <= 8'h7a;
         6311: data_out <= 8'h88;
         6312: data_out <= 8'h02;
         6313: data_out <= 8'h6e;
         6314: data_out <= 8'h7c;
         6315: data_out <= 8'h2a;
         6316: data_out <= 8'ha0;
         6317: data_out <= 8'he6;
         6318: data_out <= 8'h7e;
         6319: data_out <= 8'haa;
         6320: data_out <= 8'haa;
         6321: data_out <= 8'h50;
         6322: data_out <= 8'h7f;
         6323: data_out <= 8'h7f;
         6324: data_out <= 8'hff;
         6325: data_out <= 8'hff;
         6326: data_out <= 8'h81;
         6327: data_out <= 8'h80;
         6328: data_out <= 8'h00;
         6329: data_out <= 8'h00;
         6330: data_out <= 8'h81;
         6331: data_out <= 8'h00;
         6332: data_out <= 8'h00;
         6333: data_out <= 8'h00;
         6334: data_out <= 8'hbd;
         6335: data_out <= 8'h15;
         6336: data_out <= 8'ha4;
         6337: data_out <= 8'hce;
         6338: data_out <= 8'h18;
         6339: data_out <= 8'h99;
         6340: data_out <= 8'h8d;
         6341: data_out <= 8'h3d;
         6342: data_out <= 8'h96;
         6343: data_out <= 8'haf;
         6344: data_out <= 8'h81;
         6345: data_out <= 8'h88;
         6346: data_out <= 8'h25;
         6347: data_out <= 8'h03;
         6348: data_out <= 8'h7e;
         6349: data_out <= 8'h14;
         6350: data_out <= 8'hde;
         6351: data_out <= 8'hbd;
         6352: data_out <= 8'h16;
         6353: data_out <= 8'h5a;
         6354: data_out <= 8'h96;
         6355: data_out <= 8'h58;
         6356: data_out <= 8'h8b;
         6357: data_out <= 8'h81;
         6358: data_out <= 8'h27;
         6359: data_out <= 8'hf4;
         6360: data_out <= 8'h36;
         6361: data_out <= 8'hce;
         6362: data_out <= 8'h14;
         6363: data_out <= 8'h07;
         6364: data_out <= 8'hbd;
         6365: data_out <= 8'h13;
         6366: data_out <= 8'h1a;
         6367: data_out <= 8'hbd;
         6368: data_out <= 8'h14;
         6369: data_out <= 8'h5b;
         6370: data_out <= 8'hce;
         6371: data_out <= 8'h00;
         6372: data_out <= 8'ha3;
         6373: data_out <= 8'hbd;
         6374: data_out <= 8'h13;
         6375: data_out <= 8'h0f;
         6376: data_out <= 8'h8d;
         6377: data_out <= 8'ha7;
         6378: data_out <= 8'hce;
         6379: data_out <= 8'h18;
         6380: data_out <= 8'h9d;
         6381: data_out <= 8'h8d;
         6382: data_out <= 8'h17;
         6383: data_out <= 8'h7f;
         6384: data_out <= 8'h00;
         6385: data_out <= 8'hbb;
         6386: data_out <= 8'h32;
         6387: data_out <= 8'hbd;
         6388: data_out <= 8'h14;
         6389: data_out <= 8'hc7;
         6390: data_out <= 8'h39;
         6391: data_out <= 8'hdf;
         6392: data_out <= 8'hbd;
         6393: data_out <= 8'hbd;
         6394: data_out <= 8'h15;
         6395: data_out <= 8'ha4;
         6396: data_out <= 8'h8d;
         6397: data_out <= 8'h05;
         6398: data_out <= 8'h8d;
         6399: data_out <= 8'h08;
         6400: data_out <= 8'hce;
         6401: data_out <= 8'h00;
         6402: data_out <= 8'ha3;
         6403: data_out <= 8'h7e;
         6404: data_out <= 8'h14;
         6405: data_out <= 8'h5e;
         6406: data_out <= 8'hdf;
         6407: data_out <= 8'hbd;
         6408: data_out <= 8'hbd;
         6409: data_out <= 8'h15;
         6410: data_out <= 8'h9f;
         6411: data_out <= 8'hde;
         6412: data_out <= 8'hbd;
         6413: data_out <= 8'he6;
         6414: data_out <= 8'h00;
         6415: data_out <= 8'hd7;
         6416: data_out <= 8'hb4;
         6417: data_out <= 8'h08;
         6418: data_out <= 8'hdf;
         6419: data_out <= 8'hbd;
         6420: data_out <= 8'h8d;
         6421: data_out <= 8'hed;
         6422: data_out <= 8'hde;
         6423: data_out <= 8'hbd;
         6424: data_out <= 8'h08;
         6425: data_out <= 8'h08;
         6426: data_out <= 8'h08;
         6427: data_out <= 8'h08;
         6428: data_out <= 8'hdf;
         6429: data_out <= 8'hbd;
         6430: data_out <= 8'hbd;
         6431: data_out <= 8'h13;
         6432: data_out <= 8'h1a;
         6433: data_out <= 8'hce;
         6434: data_out <= 8'h00;
         6435: data_out <= 8'ha7;
         6436: data_out <= 8'h7a;
         6437: data_out <= 8'h00;
         6438: data_out <= 8'hb4;
         6439: data_out <= 8'h26;
         6440: data_out <= 8'heb;
         6441: data_out <= 8'h39;
         6442: data_out <= 8'h98;
         6443: data_out <= 8'h35;
         6444: data_out <= 8'h44;
         6445: data_out <= 8'h7a;
         6446: data_out <= 8'h68;
         6447: data_out <= 8'h28;
         6448: data_out <= 8'hb1;
         6449: data_out <= 8'h46;
         6450: data_out <= 8'hbd;
         6451: data_out <= 8'h15;
         6452: data_out <= 8'hd9;
         6453: data_out <= 8'h17;
         6454: data_out <= 8'h2b;
         6455: data_out <= 8'h14;
         6456: data_out <= 8'hce;
         6457: data_out <= 8'h01;
         6458: data_out <= 8'h0d;
         6459: data_out <= 8'hbd;
         6460: data_out <= 8'h15;
         6461: data_out <= 8'h8e;
         6462: data_out <= 8'h4d;
         6463: data_out <= 8'h27;
         6464: data_out <= 8'he8;
         6465: data_out <= 8'hce;
         6466: data_out <= 8'h19;
         6467: data_out <= 8'h2a;
         6468: data_out <= 8'h8d;
         6469: data_out <= 8'hbd;
         6470: data_out <= 8'hce;
         6471: data_out <= 8'h19;
         6472: data_out <= 8'h2e;
         6473: data_out <= 8'hbd;
         6474: data_out <= 8'h13;
         6475: data_out <= 8'h1a;
         6476: data_out <= 8'hd6;
         6477: data_out <= 8'hb2;
         6478: data_out <= 8'h96;
         6479: data_out <= 8'hb0;
         6480: data_out <= 8'h97;
         6481: data_out <= 8'hb2;
         6482: data_out <= 8'hd7;
         6483: data_out <= 8'hb0;
         6484: data_out <= 8'h7f;
         6485: data_out <= 8'h00;
         6486: data_out <= 8'hb3;
         6487: data_out <= 8'h96;
         6488: data_out <= 8'haf;
         6489: data_out <= 8'h97;
         6490: data_out <= 8'hbc;
         6491: data_out <= 8'h86;
         6492: data_out <= 8'h80;
         6493: data_out <= 8'h97;
         6494: data_out <= 8'haf;
         6495: data_out <= 8'hbd;
         6496: data_out <= 8'h13;
         6497: data_out <= 8'h6b;
         6498: data_out <= 8'hce;
         6499: data_out <= 8'h01;
         6500: data_out <= 8'h0d;
         6501: data_out <= 8'h7e;
         6502: data_out <= 8'h15;
         6503: data_out <= 8'haa;
         6504: data_out <= 8'hce;
         6505: data_out <= 8'h19;
         6506: data_out <= 8'hd7;
         6507: data_out <= 8'hbd;
         6508: data_out <= 8'h13;
         6509: data_out <= 8'h1a;
         6510: data_out <= 8'hbd;
         6511: data_out <= 8'h15;
         6512: data_out <= 8'hcc;
         6513: data_out <= 8'hce;
         6514: data_out <= 8'h19;
         6515: data_out <= 8'hdb;
         6516: data_out <= 8'hd6;
         6517: data_out <= 8'hba;
         6518: data_out <= 8'hbd;
         6519: data_out <= 8'h15;
         6520: data_out <= 8'h0d;
         6521: data_out <= 8'hbd;
         6522: data_out <= 8'h15;
         6523: data_out <= 8'hcc;
         6524: data_out <= 8'hbd;
         6525: data_out <= 8'h16;
         6526: data_out <= 8'h5a;
         6527: data_out <= 8'h7f;
         6528: data_out <= 8'h00;
         6529: data_out <= 8'hbb;
         6530: data_out <= 8'h96;
         6531: data_out <= 8'hb6;
         6532: data_out <= 8'hd6;
         6533: data_out <= 8'haf;
         6534: data_out <= 8'hbd;
         6535: data_out <= 8'h13;
         6536: data_out <= 8'h12;
         6537: data_out <= 8'hce;
         6538: data_out <= 8'h19;
         6539: data_out <= 8'hdf;
         6540: data_out <= 8'hbd;
         6541: data_out <= 8'h13;
         6542: data_out <= 8'h0f;
         6543: data_out <= 8'h96;
         6544: data_out <= 8'hb3;
         6545: data_out <= 8'h36;
         6546: data_out <= 8'h2a;
         6547: data_out <= 8'h0a;
         6548: data_out <= 8'hbd;
         6549: data_out <= 8'h13;
         6550: data_out <= 8'h0a;
         6551: data_out <= 8'h96;
         6552: data_out <= 8'hb3;
         6553: data_out <= 8'h2b;
         6554: data_out <= 8'h06;
         6555: data_out <= 8'h73;
         6556: data_out <= 8'h00;
         6557: data_out <= 8'h60;
         6558: data_out <= 8'hbd;
         6559: data_out <= 8'h18;
         6560: data_out <= 8'h91;
         6561: data_out <= 8'hce;
         6562: data_out <= 8'h19;
         6563: data_out <= 8'hdf;
         6564: data_out <= 8'hbd;
         6565: data_out <= 8'h13;
         6566: data_out <= 8'h1a;
         6567: data_out <= 8'h32;
         6568: data_out <= 8'h4d;
         6569: data_out <= 8'h2a;
         6570: data_out <= 8'h03;
         6571: data_out <= 8'hbd;
         6572: data_out <= 8'h18;
         6573: data_out <= 8'h91;
         6574: data_out <= 8'hce;
         6575: data_out <= 8'h19;
         6576: data_out <= 8'he3;
         6577: data_out <= 8'h7e;
         6578: data_out <= 8'h18;
         6579: data_out <= 8'hf7;
         6580: data_out <= 8'hbd;
         6581: data_out <= 8'h15;
         6582: data_out <= 8'ha4;
         6583: data_out <= 8'h7f;
         6584: data_out <= 8'h00;
         6585: data_out <= 8'h60;
         6586: data_out <= 8'h8d;
         6587: data_out <= 8'hb2;
         6588: data_out <= 8'hce;
         6589: data_out <= 8'h00;
         6590: data_out <= 8'hab;
         6591: data_out <= 8'h8d;
         6592: data_out <= 8'ha4;
         6593: data_out <= 8'hce;
         6594: data_out <= 8'h00;
         6595: data_out <= 8'ha3;
         6596: data_out <= 8'hbd;
         6597: data_out <= 8'h15;
         6598: data_out <= 8'h8e;
         6599: data_out <= 8'h7f;
         6600: data_out <= 8'h00;
         6601: data_out <= 8'hb3;
         6602: data_out <= 8'h96;
         6603: data_out <= 8'h60;
         6604: data_out <= 8'h8d;
         6605: data_out <= 8'h06;
         6606: data_out <= 8'hce;
         6607: data_out <= 8'h00;
         6608: data_out <= 8'hab;
         6609: data_out <= 8'h7e;
         6610: data_out <= 8'h15;
         6611: data_out <= 8'h12;
         6612: data_out <= 8'h36;
         6613: data_out <= 8'h20;
         6614: data_out <= 8'hc7;
         6615: data_out <= 8'h81;
         6616: data_out <= 8'h49;
         6617: data_out <= 8'h0f;
         6618: data_out <= 8'hdb;
         6619: data_out <= 8'h83;
         6620: data_out <= 8'h49;
         6621: data_out <= 8'h0f;
         6622: data_out <= 8'hdb;
         6623: data_out <= 8'h7f;
         6624: data_out <= 8'h00;
         6625: data_out <= 8'h00;
         6626: data_out <= 8'h00;
         6627: data_out <= 8'h04;
         6628: data_out <= 8'h86;
         6629: data_out <= 8'h1e;
         6630: data_out <= 8'hd7;
         6631: data_out <= 8'hba;
         6632: data_out <= 8'h87;
         6633: data_out <= 8'h99;
         6634: data_out <= 8'h26;
         6635: data_out <= 8'h64;
         6636: data_out <= 8'h87;
         6637: data_out <= 8'h23;
         6638: data_out <= 8'h34;
         6639: data_out <= 8'h58;
         6640: data_out <= 8'h86;
         6641: data_out <= 8'ha5;
         6642: data_out <= 8'h5d;
         6643: data_out <= 8'he0;
         6644: data_out <= 8'h83;
         6645: data_out <= 8'h49;
         6646: data_out <= 8'h0f;
         6647: data_out <= 8'hda;
         6648: data_out <= 8'h96;
         6649: data_out <= 8'hb3;
         6650: data_out <= 8'h36;
         6651: data_out <= 8'h2a;
         6652: data_out <= 8'h02;
         6653: data_out <= 8'h8d;
         6654: data_out <= 8'h20;
         6655: data_out <= 8'h96;
         6656: data_out <= 8'haf;
         6657: data_out <= 8'h36;
         6658: data_out <= 8'h81;
         6659: data_out <= 8'h81;
         6660: data_out <= 8'h25;
         6661: data_out <= 8'h05;
         6662: data_out <= 8'hce;
         6663: data_out <= 8'h14;
         6664: data_out <= 8'h07;
         6665: data_out <= 8'h8d;
         6666: data_out <= 8'hc6;
         6667: data_out <= 8'hce;
         6668: data_out <= 8'h1a;
         6669: data_out <= 8'h23;
         6670: data_out <= 8'h8d;
         6671: data_out <= 8'ha1;
         6672: data_out <= 8'h32;
         6673: data_out <= 8'h81;
         6674: data_out <= 8'h81;
         6675: data_out <= 8'h25;
         6676: data_out <= 8'h06;
         6677: data_out <= 8'hce;
         6678: data_out <= 8'h19;
         6679: data_out <= 8'hd7;
         6680: data_out <= 8'hbd;
         6681: data_out <= 8'h13;
         6682: data_out <= 8'h0f;
         6683: data_out <= 8'h32;
         6684: data_out <= 8'h4d;
         6685: data_out <= 8'h2a;
         6686: data_out <= 8'h03;
         6687: data_out <= 8'h7e;
         6688: data_out <= 8'h18;
         6689: data_out <= 8'h91;
         6690: data_out <= 8'h39;
         6691: data_out <= 8'h08;
         6692: data_out <= 8'h78;
         6693: data_out <= 8'h3b;
         6694: data_out <= 8'hd7;
         6695: data_out <= 8'h4a;
         6696: data_out <= 8'h7b;
         6697: data_out <= 8'h84;
         6698: data_out <= 8'h6e;
         6699: data_out <= 8'h02;
         6700: data_out <= 8'h7c;
         6701: data_out <= 8'h2f;
         6702: data_out <= 8'hc1;
         6703: data_out <= 8'hfe;
         6704: data_out <= 8'h7d;
         6705: data_out <= 8'h9a;
         6706: data_out <= 8'h31;
         6707: data_out <= 8'h74;
         6708: data_out <= 8'h7d;
         6709: data_out <= 8'h5a;
         6710: data_out <= 8'h3d;
         6711: data_out <= 8'h84;
         6712: data_out <= 8'h7e;
         6713: data_out <= 8'h91;
         6714: data_out <= 8'h7f;
         6715: data_out <= 8'hc8;
         6716: data_out <= 8'h7e;
         6717: data_out <= 8'h4c;
         6718: data_out <= 8'hbb;
         6719: data_out <= 8'he4;
         6720: data_out <= 8'h7f;
         6721: data_out <= 8'haa;
         6722: data_out <= 8'haa;
         6723: data_out <= 8'h6c;
         6724: data_out <= 8'h81;
         6725: data_out <= 8'h00;
         6726: data_out <= 8'h00;
         6727: data_out <= 8'h00;
         6728: data_out <= 8'h00;
         6729: data_out <= 8'hce;
         6730: data_out <= 8'h1b;
         6731: data_out <= 8'h75;
         6732: data_out <= 8'hbd;
         6733: data_out <= 8'h08;
         6734: data_out <= 8'h87;
         6735: data_out <= 8'hce;
         6736: data_out <= 8'hff;
         6737: data_out <= 8'hff;
         6738: data_out <= 8'hdf;
         6739: data_out <= 8'h8a;
         6740: data_out <= 8'h8e;
         6741: data_out <= 8'h1c;
         6742: data_out <= 8'h7c;
         6743: data_out <= 8'h9f;
         6744: data_out <= 8'h82;
         6745: data_out <= 8'h7f;
         6746: data_out <= 8'h01;
         6747: data_out <= 8'h11;
         6748: data_out <= 8'hbd;
         6749: data_out <= 8'h08;
         6750: data_out <= 8'h42;
         6751: data_out <= 8'hce;
         6752: data_out <= 8'h00;
         6753: data_out <= 8'h65;
         6754: data_out <= 8'hdf;
         6755: data_out <= 8'h61;
         6756: data_out <= 8'hce;
         6757: data_out <= 8'h1c;
         6758: data_out <= 8'h0b;
         6759: data_out <= 8'hbd;
         6760: data_out <= 8'h08;
         6761: data_out <= 8'h87;
         6762: data_out <= 8'hbd;
         6763: data_out <= 8'h09;
         6764: data_out <= 8'h07;
         6765: data_out <= 8'hdf;
         6766: data_out <= 8'hc8;
         6767: data_out <= 8'hbd;
         6768: data_out <= 8'h00;
         6769: data_out <= 8'hbf;
         6770: data_out <= 8'h81;
         6771: data_out <= 8'h41;
         6772: data_out <= 8'h27;
         6773: data_out <= 8'hd3;
         6774: data_out <= 8'h4d;
         6775: data_out <= 8'h26;
         6776: data_out <= 8'h15;
         6777: data_out <= 8'hce;
         6778: data_out <= 8'h1c;
         6779: data_out <= 8'h18;
         6780: data_out <= 8'h08;
         6781: data_out <= 8'h86;
         6782: data_out <= 8'h37;
         6783: data_out <= 8'ha7;
         6784: data_out <= 8'h00;
         6785: data_out <= 8'ha1;
         6786: data_out <= 8'h00;
         6787: data_out <= 8'h26;
         6788: data_out <= 8'h17;
         6789: data_out <= 8'h4a;
         6790: data_out <= 8'ha7;
         6791: data_out <= 8'h00;
         6792: data_out <= 8'ha1;
         6793: data_out <= 8'h00;
         6794: data_out <= 8'h27;
         6795: data_out <= 8'hf0;
         6796: data_out <= 8'h20;
         6797: data_out <= 8'h0e;
         6798: data_out <= 8'hbd;
         6799: data_out <= 8'h00;
         6800: data_out <= 8'hc7;
         6801: data_out <= 8'hbd;
         6802: data_out <= 8'h07;
         6803: data_out <= 8'h75;
         6804: data_out <= 8'h4d;
         6805: data_out <= 8'h27;
         6806: data_out <= 8'h03;
         6807: data_out <= 8'h7e;
         6808: data_out <= 8'h0b;
         6809: data_out <= 8'h57;
         6810: data_out <= 8'hde;
         6811: data_out <= 8'h8e;
         6812: data_out <= 8'h09;
         6813: data_out <= 8'hdf;
         6814: data_out <= 8'h88;
         6815: data_out <= 8'hdf;
         6816: data_out <= 8'h84;
         6817: data_out <= 8'hce;
         6818: data_out <= 8'h1b;
         6819: data_out <= 8'h99;
         6820: data_out <= 8'hbd;
         6821: data_out <= 8'h08;
         6822: data_out <= 8'h87;
         6823: data_out <= 8'hbd;
         6824: data_out <= 8'h09;
         6825: data_out <= 8'h07;
         6826: data_out <= 8'hdf;
         6827: data_out <= 8'hc8;
         6828: data_out <= 8'hbd;
         6829: data_out <= 8'h00;
         6830: data_out <= 8'hbf;
         6831: data_out <= 8'h16;
         6832: data_out <= 8'h27;
         6833: data_out <= 8'h1c;
         6834: data_out <= 8'hbd;
         6835: data_out <= 8'h07;
         6836: data_out <= 8'h75;
         6837: data_out <= 8'h96;
         6838: data_out <= 8'h8e;
         6839: data_out <= 8'h26;
         6840: data_out <= 8'he8;
         6841: data_out <= 8'h96;
         6842: data_out <= 8'h8f;
         6843: data_out <= 8'h81;
         6844: data_out <= 8'h10;
         6845: data_out <= 8'h25;
         6846: data_out <= 8'he2;
         6847: data_out <= 8'h97;
         6848: data_out <= 8'h0c;
         6849: data_out <= 8'h80;
         6850: data_out <= 8'h0e;
         6851: data_out <= 8'h24;
         6852: data_out <= 8'hfc;
         6853: data_out <= 8'h40;
         6854: data_out <= 8'h80;
         6855: data_out <= 8'h0e;
         6856: data_out <= 8'h9b;
         6857: data_out <= 8'h0c;
         6858: data_out <= 8'h97;
         6859: data_out <= 8'h0d;
         6860: data_out <= 8'h20;
         6861: data_out <= 8'h08;
         6862: data_out <= 8'h86;
         6863: data_out <= 8'h48;
         6864: data_out <= 8'h97;
         6865: data_out <= 8'h0c;
         6866: data_out <= 8'h86;
         6867: data_out <= 8'h38;
         6868: data_out <= 8'h97;
         6869: data_out <= 8'h0d;
         6870: data_out <= 8'hc6;
         6871: data_out <= 8'hce;
         6872: data_out <= 8'h86;
         6873: data_out <= 8'hff;
         6874: data_out <= 8'hdb;
         6875: data_out <= 8'h89;
         6876: data_out <= 8'h99;
         6877: data_out <= 8'h88;
         6878: data_out <= 8'h25;
         6879: data_out <= 8'h03;
         6880: data_out <= 8'h7e;
         6881: data_out <= 8'h03;
         6882: data_out <= 8'h1f;
         6883: data_out <= 8'h97;
         6884: data_out <= 8'h82;
         6885: data_out <= 8'hd7;
         6886: data_out <= 8'h83;
         6887: data_out <= 8'hce;
         6888: data_out <= 8'h1b;
         6889: data_out <= 8'h60;
         6890: data_out <= 8'hbd;
         6891: data_out <= 8'h08;
         6892: data_out <= 8'h87;
         6893: data_out <= 8'hbd;
         6894: data_out <= 8'h09;
         6895: data_out <= 8'h07;
         6896: data_out <= 8'hdf;
         6897: data_out <= 8'hc8;
         6898: data_out <= 8'hbd;
         6899: data_out <= 8'h00;
         6900: data_out <= 8'hbf;
         6901: data_out <= 8'hce;
         6902: data_out <= 8'h1a;
         6903: data_out <= 8'h48;
         6904: data_out <= 8'h81;
         6905: data_out <= 8'h59;
         6906: data_out <= 8'h27;
         6907: data_out <= 8'h24;
         6908: data_out <= 8'h81;
         6909: data_out <= 8'h41;
         6910: data_out <= 8'h27;
         6911: data_out <= 8'h04;
         6912: data_out <= 8'h81;
         6913: data_out <= 8'h4e;
         6914: data_out <= 8'h26;
         6915: data_out <= 8'he3;
         6916: data_out <= 8'hce;
         6917: data_out <= 8'h0d;
         6918: data_out <= 8'h71;
         6919: data_out <= 8'hff;
         6920: data_out <= 8'h01;
         6921: data_out <= 8'h33;
         6922: data_out <= 8'hce;
         6923: data_out <= 8'h19;
         6924: data_out <= 8'hf8;
         6925: data_out <= 8'h81;
         6926: data_out <= 8'h41;
         6927: data_out <= 8'h27;
         6928: data_out <= 8'h0f;
         6929: data_out <= 8'hce;
         6930: data_out <= 8'h0d;
         6931: data_out <= 8'h71;
         6932: data_out <= 8'hff;
         6933: data_out <= 8'h01;
         6934: data_out <= 8'h2d;
         6935: data_out <= 8'hff;
         6936: data_out <= 8'h01;
         6937: data_out <= 8'h31;
         6938: data_out <= 8'hff;
         6939: data_out <= 8'h01;
         6940: data_out <= 8'h2f;
         6941: data_out <= 8'hce;
         6942: data_out <= 8'h19;
         6943: data_out <= 8'h68;
         6944: data_out <= 8'h4f;
         6945: data_out <= 8'ha7;
         6946: data_out <= 8'h00;
         6947: data_out <= 8'h08;
         6948: data_out <= 8'hdf;
         6949: data_out <= 8'h7a;
         6950: data_out <= 8'hde;
         6951: data_out <= 8'h82;
         6952: data_out <= 8'h2b;
         6953: data_out <= 8'h05;
         6954: data_out <= 8'h8c;
         6955: data_out <= 8'h1c;
         6956: data_out <= 8'h7c;
         6957: data_out <= 8'h2b;
         6958: data_out <= 8'hb1;
         6959: data_out <= 8'hdf;
         6960: data_out <= 8'h82;
         6961: data_out <= 8'h96;
         6962: data_out <= 8'h7a;
         6963: data_out <= 8'hd6;
         6964: data_out <= 8'h7b;
         6965: data_out <= 8'hbd;
         6966: data_out <= 8'h02;
         6967: data_out <= 8'hfe;
         6968: data_out <= 8'hbd;
         6969: data_out <= 8'h08;
         6970: data_out <= 8'h42;
         6971: data_out <= 8'hd6;
         6972: data_out <= 8'h83;
         6973: data_out <= 8'hd0;
         6974: data_out <= 8'h7b;
         6975: data_out <= 8'h96;
         6976: data_out <= 8'h82;
         6977: data_out <= 8'h92;
         6978: data_out <= 8'h7a;
         6979: data_out <= 8'hbd;
         6980: data_out <= 8'h17;
         6981: data_out <= 8'h36;
         6982: data_out <= 8'hce;
         6983: data_out <= 8'h1b;
         6984: data_out <= 8'ha8;
         6985: data_out <= 8'hbd;
         6986: data_out <= 8'h08;
         6987: data_out <= 8'h87;
         6988: data_out <= 8'hce;
         6989: data_out <= 8'h08;
         6990: data_out <= 8'h87;
         6991: data_out <= 8'hff;
         6992: data_out <= 8'h01;
         6993: data_out <= 8'h13;
         6994: data_out <= 8'hbd;
         6995: data_out <= 8'h04;
         6996: data_out <= 8'hf2;
         6997: data_out <= 8'h86;
         6998: data_out <= 8'hbd;
         6999: data_out <= 8'h97;
         7000: data_out <= 8'h04;
         7001: data_out <= 8'hce;
         7002: data_out <= 8'h05;
         7003: data_out <= 8'h0e;
         7004: data_out <= 8'hdf;
         7005: data_out <= 8'h05;
         7006: data_out <= 8'h7e;
         7007: data_out <= 8'h03;
         7008: data_out <= 8'h4a;
         7009: data_out <= 8'h57;
         7010: data_out <= 8'h41;
         7011: data_out <= 8'h4e;
         7012: data_out <= 8'h54;
         7013: data_out <= 8'h20;
         7014: data_out <= 8'h53;
         7015: data_out <= 8'h49;
         7016: data_out <= 8'h4e;
         7017: data_out <= 8'h2d;
         7018: data_out <= 8'h43;
         7019: data_out <= 8'h4f;
         7020: data_out <= 8'h53;
         7021: data_out <= 8'h2d;
         7022: data_out <= 8'h54;
         7023: data_out <= 8'h41;
         7024: data_out <= 8'h4e;
         7025: data_out <= 8'h2d;
         7026: data_out <= 8'h41;
         7027: data_out <= 8'h54;
         7028: data_out <= 8'hce;
         7029: data_out <= 8'h00;
         7030: data_out <= 8'h0d;
         7031: data_out <= 8'h0a;
         7032: data_out <= 8'h0c;
         7033: data_out <= 8'h57;
         7034: data_out <= 8'h52;
         7035: data_out <= 8'h49;
         7036: data_out <= 8'h54;
         7037: data_out <= 8'h54;
         7038: data_out <= 8'h45;
         7039: data_out <= 8'h4e;
         7040: data_out <= 8'h20;
         7041: data_out <= 8'h42;
         7042: data_out <= 8'h59;
         7043: data_out <= 8'h20;
         7044: data_out <= 8'h52;
         7045: data_out <= 8'h49;
         7046: data_out <= 8'h43;
         7047: data_out <= 8'h48;
         7048: data_out <= 8'h41;
         7049: data_out <= 8'h52;
         7050: data_out <= 8'h44;
         7051: data_out <= 8'h20;
         7052: data_out <= 8'h57;
         7053: data_out <= 8'h2e;
         7054: data_out <= 8'h20;
         7055: data_out <= 8'h57;
         7056: data_out <= 8'h45;
         7057: data_out <= 8'h49;
         7058: data_out <= 8'h4c;
         7059: data_out <= 8'h41;
         7060: data_out <= 8'h4e;
         7061: data_out <= 8'h44;
         7062: data_out <= 8'hae;
         7063: data_out <= 8'h0d;
         7064: data_out <= 8'h0a;
         7065: data_out <= 8'h00;
         7066: data_out <= 8'h54;
         7067: data_out <= 8'h45;
         7068: data_out <= 8'h52;
         7069: data_out <= 8'h4d;
         7070: data_out <= 8'h49;
         7071: data_out <= 8'h4e;
         7072: data_out <= 8'h41;
         7073: data_out <= 8'h4c;
         7074: data_out <= 8'h20;
         7075: data_out <= 8'h57;
         7076: data_out <= 8'h49;
         7077: data_out <= 8'h44;
         7078: data_out <= 8'h54;
         7079: data_out <= 8'hc8;
         7080: data_out <= 8'h00;
         7081: data_out <= 8'h20;
         7082: data_out <= 8'h42;
         7083: data_out <= 8'h59;
         7084: data_out <= 8'h54;
         7085: data_out <= 8'h45;
         7086: data_out <= 8'h53;
         7087: data_out <= 8'h20;
         7088: data_out <= 8'h46;
         7089: data_out <= 8'h52;
         7090: data_out <= 8'h45;
         7091: data_out <= 8'hc5;
         7092: data_out <= 8'h0d;
         7093: data_out <= 8'h0a;
         7094: data_out <= 8'h0d;
         7095: data_out <= 8'h0a;
         7096: data_out <= 8'h4d;
         7097: data_out <= 8'h49;
         7098: data_out <= 8'h54;
         7099: data_out <= 8'h53;
         7100: data_out <= 8'h20;
         7101: data_out <= 8'h41;
         7102: data_out <= 8'h4c;
         7103: data_out <= 8'h54;
         7104: data_out <= 8'h41;
         7105: data_out <= 8'h49;
         7106: data_out <= 8'h52;
         7107: data_out <= 8'h20;
         7108: data_out <= 8'h36;
         7109: data_out <= 8'h38;
         7110: data_out <= 8'h30;
         7111: data_out <= 8'h20;
         7112: data_out <= 8'h42;
         7113: data_out <= 8'h41;
         7114: data_out <= 8'h53;
         7115: data_out <= 8'h49;
         7116: data_out <= 8'h43;
         7117: data_out <= 8'h20;
         7118: data_out <= 8'h56;
         7119: data_out <= 8'h45;
         7120: data_out <= 8'h52;
         7121: data_out <= 8'h53;
         7122: data_out <= 8'h49;
         7123: data_out <= 8'h4f;
         7124: data_out <= 8'h4e;
         7125: data_out <= 8'h20;
         7126: data_out <= 8'h31;
         7127: data_out <= 8'h2e;
         7128: data_out <= 8'h31;
         7129: data_out <= 8'h20;
         7130: data_out <= 8'h52;
         7131: data_out <= 8'h45;
         7132: data_out <= 8'h56;
         7133: data_out <= 8'h20;
         7134: data_out <= 8'h33;
         7135: data_out <= 8'h2e;
         7136: data_out <= 8'hb2;
         7137: data_out <= 8'h0d;
         7138: data_out <= 8'h0a;
         7139: data_out <= 8'h2d;
         7140: data_out <= 8'h2d;
         7141: data_out <= 8'h4b;
         7142: data_out <= 8'h43;
         7143: data_out <= 8'h41;
         7144: data_out <= 8'h43;
         7145: data_out <= 8'h52;
         7146: data_out <= 8'h2d;
         7147: data_out <= 8'had;
         7148: data_out <= 8'h0d;
         7149: data_out <= 8'h0a;
         7150: data_out <= 8'h43;
         7151: data_out <= 8'h4f;
         7152: data_out <= 8'h50;
         7153: data_out <= 8'h59;
         7154: data_out <= 8'h52;
         7155: data_out <= 8'h49;
         7156: data_out <= 8'h47;
         7157: data_out <= 8'h48;
         7158: data_out <= 8'h54;
         7159: data_out <= 8'h20;
         7160: data_out <= 8'h31;
         7161: data_out <= 8'h39;
         7162: data_out <= 8'h37;
         7163: data_out <= 8'h36;
         7164: data_out <= 8'h20;
         7165: data_out <= 8'h42;
         7166: data_out <= 8'h59;
         7167: data_out <= 8'h20;
         7168: data_out <= 8'h4d;
         7169: data_out <= 8'h49;
         7170: data_out <= 8'h54;
         7171: data_out <= 8'h53;
         7172: data_out <= 8'h20;
         7173: data_out <= 8'h49;
         7174: data_out <= 8'h4e;
         7175: data_out <= 8'h43;
         7176: data_out <= 8'hae;
         7177: data_out <= 8'h0d;
         7178: data_out <= 8'h0a;
         7179: data_out <= 8'h00;
         7180: data_out <= 8'h4d;
         7181: data_out <= 8'h45;
         7182: data_out <= 8'h4d;
         7183: data_out <= 8'h4f;
         7184: data_out <= 8'h52;
         7185: data_out <= 8'h59;
         7186: data_out <= 8'h20;
         7187: data_out <= 8'h53;
         7188: data_out <= 8'h49;
         7189: data_out <= 8'h5a;
         7190: data_out <= 8'hc5;
         7191: data_out <= 8'h00;
         7192: data_out <= 8'h00;
         default: data_out <= 8'h00;
      endcase
   end

endmodule

